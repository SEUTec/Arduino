    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz    ��  CPart    �����   �  �  �����   �  �              voltage_source��  CIntPin    ��  CWire   	 �        �
   /   �   �      /   �   �                  Marker ��  CExtPin    ��  CVertexA   �  �   ��  CSegment=    �G   �  �                 �:    �O   �  �   �    �"   �  �                           
        `      M     @  `          Ctrl     ��   CPin                   ��                                                           `   M��  TLine     P       `     ��    ��                                                ��  TPolygon     ����    ����   ��                                                         ��  TPoint    0        �   @        �    P        �0   @            ��  
 TTextField    �����        ��                                                          �����         �����      	[refname]       X  Q  �  �        �   ,                Marker     Miscellaneous      �?    +   ��   CMarkerBehavior     ��  CValue             0.0      �������� M ��  	 TModelPin ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      "   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               & Analog MiscV   Generic   CtrlCtrl          ����               Ctrl  v(Ctrl)  N ��   CPartPin    ����MM       A    ����RootmarkerGeneric              Ctrl �        �   /   �   �      /   �   �                  Marker) 	�    �    �  �   �/   , �   �  �   -                       `      MȘ� `  `          Ctrl     �                   ��                                                           `   M�     P       `     ��                                                        �     ����    ����   ��                                                         �    0        �   @        �    P        �0   @            �    �����        ��                                                          �����         �����      	[refname]       x  Q    �        �   ,    1   / 6 0      Marker     Miscellaneous      �?    +   !�     #�             0.0      �������� M %� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      7   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               9 Analog MiscV   Generic   CtrlCtrl          ����               Ctrl  v(Ctrl)  N '�    ����MM       A  �����RootmarkerGeneric              Ctrl �        �   /   �   �      /   �   �                  Marker; 	�    �   �  �   �   > �   �  �   ?                       `      M����    `          Ctrl     �                   ��                                                           `   M�     P       `     ��     �                                                 �     ����    ����   ��                                                         �    0        �   @        �    P        �0   @            �    �����        ��                                                          �����         �����      	[refname]       8  Q  �  �        �   ,    C   A H B      Marker     Miscellaneous      �?    +   !�     #�             0.0      �������� M %� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      I   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               K Analog MiscV   Generic   CtrlCtrl          ����               Ctrl  v(Ctrl)  N '�    ����MM       A �������RootmarkerGeneric              Ctrl �        �   /   �   �      /   �   �                  MarkerM 	�    �
   �  �   �   P �!   �  @   Q                       `      Mhz� `  �          Ctrl     �                   ��                                                           `   M�     P       `     ��                                                        �     ����    ����   ��                                                         �    0        �   @        �    P        �0   @            �    �����        ��                                                          �����         �����      	[refname]       x  �    Q        �   ,    U   S Z T      Marker     Miscellaneous      �?    +   !�     #�             0.0      �������� M %� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      [   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               ] Analog MiscV   Generic   CtrlCtrl          ����               Ctrl  v(Ctrl)  N '�    ����MM       A pH�����RootmarkerGeneric              Ctrl �      �       �   �  �      �   �  �              vcswitch�    �     �    b     �           �   �           �   �               Gndc 	�    �H   @  �   �   �I   @  `   g         f     �   �J      �   �8   �      �
   k         j     �#   �D   �   �   �5   �   �   `	   o         n     m      j     i      f     �   f �4    
  �   �   �L    
  `   s          r     q �   r �9      �   �   �      `   w          v     u �   v �1      �   �   �M      �   �   �N      `   }      |     {          z     y                                        `       Gnd}   �  �          gnd1     �                    ��                                                               Gnd�                   ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��    p�Z         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ          � � �   �      Ground    
Ground DINMiscellaneous      �?       ��   CGroundBehavior       Gnd ��   CBehPin     Gnd        ����Gnd����                        ��gndgnd                 � Analog Meters   Generic   gnd1gnd1          ����  gnd '�    ����GndGnd      GNDAGnd �)����SourcesGroundGeneric              0 �   b    �       �   �  �      �   �  �              vcswitch�    �    �    �   �       _   �         _   �                 capacitor_generic� �   �    � �   �   �       S   �  ,      S   �  ,              Ammeter�    �    �   �   �       �   �        �   �                Inductor�    �    �    �    �       �   �  �       �   �  �               R� �   �   � 3 	�    �   �
  @   �-   � �      @   �                        �  �   R+  	�   �   `	  @   �,   �7   @  @   � �7   �=   @  �	   �3   � �8   �
  �	   �            � �   �5   @  @   �$   � �      @   �             �%   �'   @  �   �;   � �&    
  �   � �   �+    
  @   �         �             �)   �>   @  `   �         �     �     �     �     �         �     �   � �3   @  `   �9   � �2    
  `   � �   � �F    
  @   �                    � �   � �   @  �   �                         �                  �   R-   `	  �
         R     �                    ��                                                       �   @   R+�                   ��                                                          @   R-�    @   $   0     ��    ��)                                                � 0   P   $   0     ��                                                        � 0   P   <   0     ��    ��)                                                � H   P   <   0     ��    p�Z                                                � H   P   T   0     ��                                                       � `   P   h   @     ��    D�Z                                                � �   @   h   @     ��    ��d                                                � `   P   T   0    	 ��    |�f	                                                �    @       @    
 ��    <�b
                                                � ����F   X   f     ��                                                       ����F   X   f   ����F   X   f   [resistance]       �  R  �	  �      `   �   �   �         t   $     ��                                                               t   $           t   $   	[refname]       `	  �
  �	             t   $    � � � � � � � � � � � � �    resistor    resistor DINMiscellaneous      �?       ��  CResistorBehavior     #� �������(\��?0.58      ��������#� ���� 27     ��������#� ����       ��������#� ����       �������� R+R- ��     R+        ����R+����                        ����    R-      ����R-����                        �� resistor                � � Passive   Generic   RR          ����    R '�    ����R+R+      PASAR+JV1.����'�   ����R-R-      PASAR-�)����Passivedefault resistor, 1KGeneric              5 �  � ��     L+        ����L+����                        �� 5   � 5 � 	�    �        �   L+K  	�   �   �  @   �.   � �.   �  @   �                      �  �   L-L      �
          L1     �                    ��                                                           @   L+�                   ��                                                      �   @   L-��   TArc h   ,   �   T    
                                                           h   ,   �   T   h   ,   �   T   �   @   h   @           ۀ P   ,   h   T    	                                                           P   ,   h   T   P   ,   h   T   h   @   P   @           ۀ 8   ,   P   T                                                               8   ,   P   T   8   ,   P   T   P   @   8   @           ۀ     ,   8   T                                                                   ,   8   T       ,   8   T   8   @       @           � $   P      X     ��    ��                                                �    H   $   P     ��     �                                                  �     P   $   P     ��    ��                                                �     @       @     ��    p�H	                                                � �   @   �   @     ��       
                                                �     \   �   |     ��                                                           \   �   |       \   �   |   [Inductance]          �  �  *      \   �   |   �         �   $     ��                                                               �   $           �   $   	[refname]          �
  p             �   $    � � �   �   �   �   � � �   �   �   �   �      Inductor     Miscellaneous      �?    
   ��  CInductorBehavior     #� ��� {�G�zt?5m      ��������#� ���� x     �������� L+L- � ��    L-      ����L-����                        �� Inductor  
              � � Passive   Generic   L1L1          ����  L '�    ����L+L+      PASAL+�4T����'�   ����L-L-      PASAL-������PassiveInductorGeneric              11 �  � ��     M+        ����M+����                        �� 11   � 11 � 	�    �        �   M+0  	�   �   @  @   �1   � �;      @   � �   �<      �	   �!   �%   �  �	   �         �     � �   �@      @   �   �-   �  @   �        �     �   �/      �   �4   �:   �  �   � �'   �C   �  @            �         �     �    �	      `          �     �     �     �     �         �     �
   � �,      `   �   �)      @              �   �K      `   �"   	�      @   
                                            �  �   M-1   �  �
          VA_IL    	 �                   ��                                                           @   M+�                   ��                                                      �   @   M-� �   @   �   @     ��    ��                                                �     @       @     ��                                                        � 4   X   `   X     ��    ��                                                �� 
 TRectangle        �   d                   ����                                                �   d   � ����������������  ��          @ @                                           �d   X    IX1.�X   P        �X   `    0000@ @ � $   $   �   L     ��                                                      $   $   �   L   $   $   �   L   [value]         �
  �  �  $   $   �   L   �     �����        ��                                                           �����          �����      	[refname]          \
    �
      �����               	     Ammeter    Ammeter_smallMiscellaneous      �?       ��   CAmmeterBehavior     #� ����   @?��-1.52      �������� M+M- � ��    M-      ����M-����                        ��AmmeterAmmeter   �            � Analog Meters   Generic   VA_ILVA_IL          ����  VAm '�    ����M+M+      PASAM+0�M����'�   ����M-M-      PASAM- ������Analog MetersAmmeterGeneric              13 �   �   ` 13 �   �   �       �   �         �   �                 1n4007�    b     !0  	�    x        @  D+   	�            D-                 D2     �                   ��                                                           �   D+�                   ��                                                          `   D-� �����       �      ��    ���                                                 �     �       �     ��                                                        � �����       �     ��    ���                                                 �     �       �     ��    (�K                                                � �����       �     ��                                                       �     �      �     ��    ��K                                                �     �       `     ��    ��K                                                � d   �   $  �    	 ��        	                                               0   `   �   �   0   `   �   �   	[devname]        �������������������������      � 0   �   �   �    
 ��        
                                               0   �   �   �   0   �   �   �   	[refname]       �  �  0  |  ����   �   <    '()*+,-    ./          %& �
  diode     Miscellaneous      �?       ��  CDiodeBehavior     #� ����  F      ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     �������� D+D- ��     D+        ����D+����                        ����    D-      ����D-����                        ��d1n4007d1n4007   S          67Diode   Generic   D2D2                D '�    ����D+D+      PASAAPKT����'�   ����D-D-      PASAK�)�����DiodeDiode	FairchildDO-41             13 �   �   �       �   �  �      �   �  �              	voltmeter�    �    ;3 :	�    �           M+i  	�   �   �     M-j                 IV_VL    
 �                   ��                                                           `   M+�                   ��                                                      �   `   M-�     `       `     ��    ��                                                � �   `   �   `     ��                                                        �    L      \     ��    ��                                                �     T      T     ��    p�H                                                � �   X   �   X     ��               	FIXED_ROT                                        �     <   �   �                   ����                                             <   �   �   � (   D   �   x     ��                                                      (   D   �   x   (   D   �   x   [value]       x  �  �  �  (   D   �   x   �        �   0    	 ��        	                                                      �   0          �   0   	[refname]       `  D  x  �         �   0    F  ?@AGC  DHE      B
     	voltmeter    voltmeter_smallMiscellaneous      �?       ��   CVoltmeterBehavior     #� �        �>476.84n      �������� M+M- ��     M+        ����M+����                        ����    M-      ����M-����                        ��	voltmeter	voltmeter   _            LMAnalog Meters   Generic   IV_VLIV_VL          ����  IVm '�    ����M+M+      PASAM+    ����'�   ����M-M-      PASAM-    ����Analog Meters Generic              13 �    �    �       �   �         �   �                 1n4007P�   �    �   S  �       _   @  �      _   @  �              Ammeter2�    �    �    W   �           �   �          �   �              BatteryX�   b    Y0 	�    �      `	   �+   �      �   ]        \               `       1�  	�   l   `   �  2�   �  `	          XSource     �                    ��                                                               1�                   ��                                                          �   2�             $     ��    ��)                                                �     \       �     ��                                                        �    8   0   8    	 ��    ��)                                                �     H   @   H     ��    p�Z                                                �     $   @   $     ��                                                       �    \   0   \     ��    D�Z                                                �               ���                                                      �               ���   �Z	                                                � `          $    
 ��        
                                               `          $   `          $   	[devname]        ����������������`          $   � `   $      H     ��                                                       `   $      H   `   $      H   	[refname]       �  �	  `  l
  `   $      H    `abcfghi    jk    e  d     Battery     Miscellaneous      �?    9 
 ��  CParamSubBehavior     #� ����      (@12      �������� 12 ��     1       ����1����                        ����    2      ����2����                        ��BatteryBattery
 9 i             opSources   Generic   XSourceXSource          ������   CParamSubModelType��    BATTERY2.SUBCKT Xbattery 1 2
V1 1 2 DC {voltage}
.ENDS
   ��  	 CParmDefn    1battery voltage   ParamSubvoltageV                X '�    ����11      PASA1�1b����'�   ����22      PASA20Ab����SourcesBatteryGeneric              4 V o��     M+        ����M+����                        �� 4   U4 T	�    ^   `   �  M+2  	�   �      `   �(   �6      @   {�*   �Q   �   @   �<   ~�(   �   �               }    |    �2   |�P   @  @   �   ��#   @  �   �           ��	   ��$    
  @   �&   ��*    
      �           ��   ��?   �  @   �0   ��B   �      �           ��   ��E      @   �6   ��      �   �            �                                    z             `   `   M-3   �            VA_Ix1    	 �                    ��                                                           �   M+�                   ��                                                              M-�     �       �     ��                                                        �     <             ��                                                        � @   <   �����                  ����                                         ����<   @   �   � ����x   ����L     ��                                                        �  ������� �������  ��          @ @                                           �����H    ��b�����T    
>DA�����T    uT@ @ � ����D   <   |     ��                                                      ����D   <   |   ����D   <   |   [value]       �  �    b     D   �   |   � ��������O        ��                                                       ��������O      ��������O      	[refname]       m  �  �       �����      
 ������  ���	   Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       �     #�  ֤�   �œC�-597.45u      �������� M+M- w��    M-      ����M-����                        ��AmmeterAmmeter   V            w�Analog Meters   Generic   VA_Ix1VA_Ix1          ����  VAm '�    ����M+M+      PASAM+��W����'�   ����M-M-      PASAM-8�W����Analog MetersAmmeter-verticalGeneric              9 �    S   �       _   �  �      _   �  �              
Voltmeter2��   b    �0 	�    �   `   `   M+k  	�   p   `   �  M-l   `   �          IV_Vx1    
 �                    ��                                                               M+�                   ��                                                          �   M-�     �       �     ��    ��                                                �             <     ��    
NVA                                                �    $      4     ��    ��                                                �    ,      ,     ��    p�H                                                �    �      �     ��               	FIXED_ROT                                        �     <   �   �                  ����                                             <   �   �   �    D   �   x     ��                                                         D   �   x      D   �   x   [value]       l   L  d  �     D   �   x   � 8      �   0    	 ��        	                                               8      �   0   8      �   0   	[refname]         �  X  D  8      �   0    �������    �      �  �
     Voltemeter-Vert    Voltemeter-Vert_smallMiscellaneous      �?       I�     #� ����      (@12.00      �������� M+M- ��     M+        ����M+����                        ����    M-      ����M-����                        ��	voltmeter	voltmeter   k            ��Analog Meters   Generic   IV_Vx1IV_Vx1          ����  IVm '�    ����M+M+      PASAM+@������'�   ����M-M-      PASAM-�����Analog MetersVoltmeter-verticalGeneric              9 �   S  �       �   �  �      �   �  �              vcswitch�    �    �3 ��      �Ctrl �   b    �0 	�    �    �   �  1S  	�   �  �      2T  	�             3U  	�   �   �  `                       �  4V   �  �        X1     �                    ��                                                       @   �   1�                   ��                                                      @   `   2�                   ��                                                          `   3�                   ��                                                          �   4�     �       �     ��                                                        �     `       �     ��                                                        �     �       �    
 ���                                                       � �����      �    	 ���                                                       ��  TEllipse D   �   <   �                  ����                                         <   �   D   �   <   �   D   �   �    �   �����               	   ����                                         �����      �   � @   `   @   �     ��        
                                                � 0   �   @   �     ��                                                        � @   �   @   �     ��                                                        �    �   �����     ��  �             	FIXED_ROT                                        �    �   4   �     ��                                                        � `   �   �   �     ��                                                       `   �   �   �   `   �   �   �   	[refname]       �  |  	        (   t   L   �     �  <    ��                                                       `   `   �   �   `   `   �   �   	[devname]        ����������������       �   (    �������      ��  �������    � �  vcswitch     Miscellaneous      �?   9 
 l�    #� �����������?1.3      ��������#� ����333333�?1.45     ��������#� ����      �?0.5     ��������#� ����    ��.A1meg     �������� 1234 ��     1       ����1����                        ����    2      ����2����                        ����    3      ����3����                        ����    4      ����4����                        ��X6_vcswitchX6_vcswitch
 9               ����Switches   Generic   X1X1          ����q���voltage controlled switch   VCSW{.subckt vcsw 1 2 3 4
S 1 2 3 4 switch
.model switch sw (vt={(Von+Voff)/2} vh={(Von-Voff)/2} ron={Ron} roff={Roff})
.ends   s�    1turnon voltage   ParamSubVon               s�    1turnoff voltage   ParamSubVoffV             s�    0on resistance   ParamSubRonOhm             s�    0off resistance   ParamSubRoffOhm               X '�    ����11      PASA18Lk����'�   ����22      PASA2    ����'�   ����33      PASA3G1  ����'�   ����44      PASA4VA_I����Switches Generic              9 �   S  �       �   �         �   �                 1n4007�    �    �3 �	�    �        @  D+   	�   �         D-     
            D1     �                   ��                                                           �   D+�                   ��                                                          `   D-� �����       �      ��    ���                                                 �     �       �     ��                                                        � �����       �     ��    ���                                                 �     �       �     ��                                                       � �����       �     ��    ��K                                                �     �      �     ��    ��K                                                �     �       `     ��                                                        � d   �   $  �    	 ��        	                                               0   `   �   �   0   `   �   �   	[devname]        �������������������������      � 0   �   �   �    
 ��        
                                               0   �   �   �   0   �   �   �   	[refname]       �
  �  0  \  ����   �   <    �������    ��          �� �
  diode     Miscellaneous      �?       0�     #� ����  F      ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     �������� D+D- ��     D+        ����D+����                        ����    D-      ����D-����                        ��d1n4007d1n4007   S          ��Diode   Generic   D1D1                D '�    ����D+D+      PASAAh~�����'�   ����D-D-      PASAK � ����DiodeDiode	FairchildDO-41             9 R�    S   �       �   �  �      �   �  �              vcswitch��   �   �13 �   b    �0 �      �Ctrl 	�    �          1S  	�         �  2T  	�   �    �  `                   �   �  3U  	�   .   �      4V      �        X3     �                    ��                                                           `   1�                   ��                                                          �   2�                   ��                                                      @   �   3�                   ��                                                      @   `   4� @   �   @   `     ��                                                        � @   �   @   �     ��                                                        � @   �   @   �    
 ���                                                       � H   �   8   �    	 ���                                                       Ɂ �����      �                  ����                                         �����      �   �����      �   � 0   �   P   �               	   ����                                         0   �   P   �   �     �       �     ��    D�H
                                                �    �       �     ��                                                       �     �       `     ��                                                        � 8   �   H   �     ��  �             	FIXED_ROT                                        � ,   �      �     ��                                                        � `   �   �   �     ��                                                       `   �   �   �   `   �   �   �   	[refname]          |  �        (   t   L   �     �  <    ��                                                       `   `   �   �   `   `   �   �   	[devname]        ����������������       �   (    	
             �  vcswitch     Miscellaneous      �?   9 
 l�    #� ����333333�?1.45      ��������#� �����������?1.3     ��������#� ����      �?0.5     ��������#� ����    ��.A1meg     �������� 1234 ��     1       ����1����                        ����    2      ����2����                        ����    3      ����3����                        ����    4      ����4����                        ��vcswitchvcswitch
 9                !Switches   Generic   X3X3          ����q���voltage controlled switch   VCSW{.subckt vcsw 1 2 3 4
S 1 2 3 4 switch
.model switch sw (vt={(Von+Voff)/2} vh={(Von-Voff)/2} ron={Ron} roff={Roff})
.ends   s�    1turnon voltage   ParamSubVon               s�    1turnoff voltage   ParamSubVoffV             s�    0on resistance   ParamSubRonOhm             s�    0off resistance   ParamSubRoffOhm               X '�    ����11      PASA1IX1.����'�   ����22      PASA2    ����'�   ����33      PASA3U  ����'�   ����44      PASA4  � ����Switches Generic              9  ������    D-      ����D-����                        �� 9  Q9 	�           @  D+   	�   �         D-    �            D3     �                   ��                                                           �   D+�                   ��                                                          `   D-� �����       �      ��    ���                                                 �     �       �     ��                                                        � �����       �     ��    ���                                                 �     �       �     ��    (�K                                                � �����       �     ��                                                       �     �      �     ��    ��K                                                �     �       `     ��    ��K                                                � d   �   $  �    	 ��        	                                               0   `   �   �   0   `   �   �   	[devname]        �������������������������      � 0   �   �   �    
 ��        
                                               0   �   �   �   0   �   �   �   	[refname]         �  �  \  ����   �   <    0123456    78          ./ �
  diode     Miscellaneous      �?       0�     #� ����  F      ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     �������� D+D- ��     D+        ����D+����                        ��+d1n4007d1n4007    �          >+Diode   Generic   D3D3                D '�    ����D+D+      PASAA   `����'�   ����D-D-      PASAK��P����DiodeDiode	FairchildDO-41             13   ��    C-      ����C-����                        ��M7>��    2      ����2����                        �� 13   � 13 	�    �   �  �   C-�  	�   �        �   C+�   �
   	          C1     �                   ��                                                       �   @   C-�                   ��                                                          @   C+�     @   @   @      ��    ���                                                 � @       @   `     ��    �b�                                                � `       `   `     ��    ���                                                 � `   @   �   @     ��    (�K                                                �     `   �   �     ��                                                           `   �   �       `   �   �   [capacitance]       �
   
  �  �
      `   �   �   �         �   $     ��                                                               �   $           �   $   	[refname]       �
   	  `  �	          �   $    GHIJK    L      EF     	Capacitor     Miscellaneous      �?       ��  CCapacitorBehavior     #� '  �dy���=20p      ��������#� ���� x     ��������#� ����       ��������#� ����       �������� C+C- ��     C+        ����C+����                        ��A 	capacitor                SAPassive   Generic   C1C1          ����  C '�    ����C+C+      PASAC+�R����'�   ����C-C-      PASAC-P�����Passive Generic              3 � �   �   �       �   �         �   �                 1n4007�    b     W0 V	�    t        @  D+   	�   �          D-     
            D4     �                   ��                                                           �   D+�                   ��                                                          `   D-� �����       �      ��    ���                                                 �     �       �     ��                                                        � �����       �     ��    ���                                                 �     �       �     ��                                                       � �����       �     ��    ��K                                                �     �      �     ��    ��K                                                �     �       `     ��                                                        � d   �   $  �    	 ��        	                                               0   `   �   �   0   `   �   �   	[devname]        �������������������������      � 0   �   �   �    
 ��        
                                               0   �   �   �   0   �   �   �   	[refname]       �
  �  0  |  ����   �   <    ]^_`abc    de          [\ �
  diode     Miscellaneous      �?       0�     #� ����  F      ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     �������� D+D- ��     D+        ����D+����                        ����    D-      ����D-����                        ��d1n4007d1n4007    @          klDiode   Generic   D4D4                D '�    ����D+D+      PASAA    ����'�   ����D-D-      PASAK    ����DiodeDiode	FairchildDO-41             3 � <�� S� L��l��     1       ����1����                        �� 3   � 3 � �   b    � 0 �      � Ctrl 	�    �    �      1S  	�   h   �   �  2T  	�   �0   �  `   �   u�   �  �   v    	                       �  3U  	�   @          4V   �  �         X4     �                    ��                                                       @   `   1�                   ��                                                      @   �   2�                   ��                                                          �   3�                   ��                                                          `   4�     �       `     ��    ���                                                 �     �       �     ��    T�W                                                �     �       �    
 ���   ���                                                 � �����      �    	 ���   (�K                                                Ɂ D   �   <   �                  ����                                         <   �   D   �   <   �   D   �   �    �   �����               	   ����                                         �����      �   � @   �   @   �     ��       
                                                � 0   �   @   �     ��    ��K                                                � @   �   @   `     ��                                                       � �����      �     ��  � ԎK        	FIXED_ROT                                        �    �   4   �     ��                                                        � T   �   �   �     ��                                                       T   �   �   �   T   �   �   �   	[refname]       |  |  �        (   t   L   � �   �   4  �     ��                                                       T   `   �   �   T   `   �   �   	[devname]        ����������������       �   (    yz{|���      ~�  �����}    � �
  vcswitch     Miscellaneous      �?   9 
 l�    #� ����333333�?1.45      ��������#� ����      �-1     ��������#� ����      �?0.5     ��������#� ����    ��.A1meg     �������� 1234 o��    2      ����2����                        ����    3      ����3����                        ����    4      ����4����                        ��X2_vcswitchX2_vcswitch
 9               o���Switches   Generic   X4X4          ����q���voltage controlled switch   VCSW{.subckt vcsw 1 2 3 4
S 1 2 3 4 switch
.model switch sw (vt={(Von+Voff)/2} vh={(Von-Voff)/2} ron={Ron} roff={Roff})
.ends   s�    1turnon voltage   ParamSubVon               s�    1turnoff voltage   ParamSubVoffV             s�    0on resistance   ParamSubRonOhm             s�    0off resistance   ParamSubRoffOhm               X '�    ����11      PASA1�>
����'�   ����22      PASA2�V�����'�   ����33      PASA3 � ����'�   ����44      PASA4 � ����Switches Generic              0 Z�X"a �    b     �           �   �           �   �               Gnd�	�       `       Gnd}   `  `          gnd2     �                    ��                                                               Gnd�                   ��    ��         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         ����  �     Ground    
Ground DINMiscellaneous      �?       ��       Gnd ��     Gnd        ����Gnd����                        ��gndgnd                 �Analog Meters   Generic   gnd2gnd2          ����  gnd '�    ����GndGnd      GNDAGnd    ����SourcesGroundGeneric              0 �    b     �	           �   �           �   �               Gnd�	�    w   `       Gnd}      �          gnd3     �                    ��                                                               Gnd�                   ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         ����  �     Ground    
Ground DINMiscellaneous      �?       ��       Gnd ��     Gnd        ����Gnd����                        ��gndgnd                 �Analog Meters   Generic   gnd3gnd3          ����  gnd '�    ����GndGnd      GNDAGnd    ����SourcesGroundGeneric              0 p�    b     �           �   �           �   �               Gnd�	�    �   �  `                     `       Gnd}   @  `          gnd4     �                    ��                                                               Gnd�                   ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��    D�H         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��    x�W         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��    X��         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         ����  �     Ground    
Ground DINMiscellaneous      �?       ��       Gnd ��     Gnd        ����Gnd����                        ��gndgnd                 �Analog Meters   Generic   gnd4gnd4          ����  gnd '�    ����GndGnd      GNDAGnd    ����SourcesGroundGeneric              0 �   b     0 �    b     �           �   �           �   �               Gnd�	�    �   `       Gnd}      `          gnd5     �                    ��                                                               Gnd�                   ��    p�H         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��    D�H         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         ����  �     Ground    
Ground DINMiscellaneous      �?       ��       Gnd ��     Gnd        ����Gnd����                        ��gndgnd                 �Analog Meters   Generic   gnd5gnd5          ����  gnd '�    ����GndGnd      GNDAGnd�����SourcesGroundGeneric              0 ��    b     �           �   �           �   �               Gnd�	�    �   �  �                    `       Gnd}   `  �          gnd6     �                    ��                                                               Gnd�                   ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��       0         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��       �         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         ����  �     Ground    
Ground DINMiscellaneous      �?       ��       Gnd ��     Gnd        ����Gnd����                        ��gndgnd                 �Analog Meters   Generic   gnd6gnd6          ����  gnd '�    ����GndGnd      GNDAGnd��������SourcesGroundGeneric              0 �   b    ` 0  ��    V-      ����V-����                        ��p� ���6����k����     1       ����1����                        ����    4      ����4����                        ��   0    ` 0 _ �	�    |        �  1S  	�            2T  	�   R   �      3U  	�   �  �   �  4V                X2     �                    ��                                                           �   1�                   ��                                                          `   2�                   ��                                                      @   `   3�                   ��                                                      @   �   4� @   �   @   �     ��    ���                                                 � @   `   @   �     ��    |-S                                                � @   �   @   �    
 ���   ���                                                 � H   �   8   �    	 ���   (�K                                                Ɂ    �   �����                  ����                                         �����      �   �����      �   � P   �   0   �               	   ����                                         0   �   P   �   �     `       �     ��       
                                                �    �       �     ��    ��K                                                �     �       �     ��                                                       � 8   �   H   �     ��  � ԎK        	FIXED_ROT                                        � ,   �      �     ��                                                        � `   �   �   �     ��                                                       `   �   �   �   `   �   �   �   	[refname]          �  �  |      (   t   L   � `   `   �   �     ��                                                       `   `   �   �   `   `   �   �   	[devname]        ����������������       �   (    �������      ��  �������    � �  vcswitch     Miscellaneous      �?   9 
 l�    #� ����333333�?1.45      ��������#� ����      �-1     ��������#� ����      �?0.5     ��������#� ����    ��.A1meg     �������� 1234 �B��    3      ����3����                        ���X5_vcswitchX5_vcswitch
 9               �B��Switches   Generic   X2X2          ����q���voltage controlled switch   VCSW{.subckt vcsw 1 2 3 4
S 1 2 3 4 switch
.model switch sw (vt={(Von+Voff)/2} vh={(Von-Voff)/2} ron={Ron} roff={Roff})
.ends   s�    1turnon voltage   ParamSubVon               s�    1turnoff voltage   ParamSubVoffV             s�    0on resistance   ParamSubRonOhm             s�    0off resistance   ParamSubRoffOhm               X '�    ����11      PASA1�� ����'�   ����22      PASA2 � ����'�   ����33      PASA3   �����'�   ����44      PASA4@
G3����Switches Generic              Ctrl q �	 ��     V+        ����V+����                        ��& 9 K �] ��! Ctrl    Ctrl �	�               V+g  	�   �      �  V-h   �  �         V1     �                   ��                                                           `   V+�                   ��                                                          �   V-Ɂ     �   �����                   ����                                         �����       �   �����       �   �    �   �����     ��    ��)                                                �     �       �     ��    ��`                                                �     �       �     ��    ��)                                                �     \       �     ��    p�Z                                                � �����   
   �    
 ��               	FIXED_ROT                                        � \   `   \   `     ��                                                      \   `   \   `   \   `   \   `           �  �  �  �                � 0   �   �   �     ��        	                                               0   �   �   �   0   �   �   �   [dc]       0  p  h            p   @   � 0   \   �   �    	 ��        
                                               0   \   �   �   0   \   �   �   	[refname]       0  �  �  t      ����t         	
            �  Voltage Source    Voltage Source DINRoot      �?       ��  CVSourceBehavior     #� ����        0      ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       �������� V+V- ��volt_sourcevolt_source   +0            ��Sources   Generic   V1V1          ����       #�0            0      ��������#�0����      @5     ��������#�0            0     ��������#�0'  ���ư>1u     ��������#�0'  ���ư>1u     ��������#�0 -1����Mb`?2m     ��������#�0 '�~j�t��?12m     ��������    #�0            0      ��������#�0����      �?1.5     ��������#�0����      I@50     ��������#�0            0     ��������#�0            0     ��������    #�0            0      ��������#�0����      �?1     ��������#�0����      �?1     ��������#�0            0     ��������#�0����      �?1     ��������    #�0            0      ��������#�0����      �?1     ��������#�0            0     ��������#�0 N  �����>2u     ��������#�0'  ���ư>1u     ��������#�0'  ���ư>1u     ��������    #�  ���� 0 0      ��������                0      �������� ����       �������� ����       �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������               V '�    ����V+V+      PWR+AV+ � ����'�   ����V-V-      PWR-AV-NDDA����Sources Generic              � Y� d ;U  �� �* <   !���N �    � � �QW� ` �   b  � � W� S� > ; >       s y �� �� Q � u ? � vg { � �i w � � } q � � � � 
m � � � {� }]� � � - �� �� � o �� k �  �  R K R l �  � .   �  P �> �  � � \  � �   ^@ � p x � wz  , R  ��� � � ��� � � � uz � � r � |� � v � � � � � ��  �n ��  f h j 	t | ~  �~             
 #�@ ����        ��������#�             0     ��������#� ����      @5     ��������#�  ʚ;�������?.1     ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true
     ��������#� ����  false     ��������               
                  #� ����        ��������#� ����       ��������#�  ����       ��������#�@ ����       ��������#�@ ����       ��������               
                  #� ����        ��������#� ����       ��������#�@ ����       ��������#�  ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������               
                 #� ����dec     ��������#� ����     @�@1k     ��������#� ����    ��.A1meg     ��������#� ����       20     ��������#� ���� true     ��������#� ���� true     ��������#� ���� true	     ��������#� ����  false
     ��������               
                 #�  ����        ��������#�  ����       ��������#�  ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������               
                  	 #� ����        ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������               
                 #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
                    #�             0      ��������#�  ��{�G�z�?40m     ��������#�  � -C��6
?0.05m     ��������#�  � -C��6
?0.05m     ��������#� ���� True     ��������#� ����  F     ��������#� ���� true     ��������#� ����  false     ��������               
                 #� ����     @�@1K      ��������#�  ����       ��������#�  ����       ��������#�  ����       ��������               
         ��              #�  ����        ��������              
                  #�  ����        ��������              
                                  
                 #�@ ����        ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true	     ��������#� ����  false
     ��������#� ���� true     ��������#� ����  false     ��������               
                 #� ����       5      ��������#� ����       5     ��������#� ����       5     ��������#� ����       5     ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#�@ ����       ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#� ���� true     ��������#� ���� true     ��������#� ����  false     ��������#� ���� true     ��������#� ����  false      ��������#� ���� true!     ��������#� ����  false"     ��������               
                        #� ����       5      ��������#� ����       5     ��������#� ����       5     ��������#� ����       5     ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#�@ ����       ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#� ���� true     ��������#� ���� true     ��������#� ����  false     ��������#� ���� true     ��������#� ����  false      ��������#� ���� true!     ��������#� ����  false"     ��������               
                 #� ����       5      ��������#� ����       5     ��������#� ����       5     ��������#� ����       5     ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#�@ ����       ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#� ���� true     ��������#� ���� true     ��������#� ����  false     ��������#� ���� true     ��������#� ����  false      ��������#� ���� true!     ��������#� ����  false"     ��������               
                 #� ����       5      ��������#� ����       5     ��������#� ����       5     ��������#� ����       5     ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#�@ ����       ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#� ���� true     ��������#� ���� true     ��������#� ����  false     ��������#� ���� true     ��������#� ����  false      ��������#� ���� true!     ��������#� ����  false"     ��������               
                 #�@ ����        ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����decade     ��������#� ���� true     ��������#� ���� true     ��������#� ���� true     ��������#� ����  false     ��������               
                 #� ����        ��������#� ����       ��������#�@ ����       ��������#�  ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������               
                        #� ����dec     ��������#� ����     @�@1k     ��������#� ����    ��.A1meg     ��������#� ����       20     ��������#� ����        0     ��������#� ����        0     ��������#� ���� true	     ��������#� ���� true
     ��������#� ����      I@50     ��������#� ���� true     ��������#� ����  false     ��������               
                         / #� ���� x'     ��������#�     �-���q=1E-12     ��������#� @B -C��6?1E-4     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x	     ��������#� ���� x!     ��������#� ����    �  500
     ��������#� ���� x     ��������#� ����    �  500     ��������#� ���� x$     ��������#� ���� x$     ��������#� ���� x%     ��������#� ���� x"     ��������#�  ���� x*     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x&     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x+     ��������#� ���� x,     ��������#� ���� x-     ��������#� ���� xg     ��������#� ���� xf     ��������#� ���� xd     ��������#� ���� xe     ��������#� ���� xh     ��������#� ���� xj     ��������#� ���� xi     ��������#� ���� xk     ��������#� ����    e��A1Gl     ��������#�             0�     ��������#� ����      @5�     ��������#� ����      @2.5�     ��������#� ����      �?.5�     ��������#� ����      @4.5�     ��������#� 
   ��&�.>1n�     ��������#� 
   ��&�.>1n�     ��������#� 
   ��&�.>1n�     ��������#� 
   ��&�.>1n�     ��������           ��  CPrimitiveModel    d1n4007   #�    1�a��%>2.55e-9      ��������#� ���� 27     ��������#�  �/�$��?0.042     ��������#� ����      �?1.75     ��������#�  �  ��v��(�>5.76e-6     ��������#�     �]}IW�=1.85e-11     ��������#� ����      �?0.75     ��������#� ����Zd;�O�?0.333     ��������#� ���� 1.11	     ��������#� ���� 3.0
     ��������#�      0     ��������#� ���� 1     ��������#� ���� 0.5     ��������#� ����     @�@1000     ��������#� � Ǯ���?9.86e-5     ��������     Diode Generic��   CPrimitiveModelType Junction Diode model����DD   s����� 1.0E-14Saturation current    ProcessisAmp0       e     s����� 27!Parameter measurement temperature    ProcesstnomDeg C0     s     s����� 0Ohmic resistance    ProcessrsOhm0      f     s����� 1Emission Coefficient    Processn 0      g     s����� 0Transit Time    Processttsec0     h     s����� 0Junction capacitance    ProcesscjoF0     i     s����� 0     Processcj0F0     i     s����� 1Junction potential    ProcessvjV0      j     s����� 0.5Grading coefficient    Processm 0      k     s����� 1.11Activation energy    ProcessegeV0     	 l     s����� 3.0#Saturation current temperature exp.    Processxti 0     
 m     s����� 0flicker noise coefficient    Processkf 0      t     s����� 1flicker noise exponent    Processaf 0      u     s����� 0.5#Forward bias junction fit parameter    Processfc 0      n     s����� infReverse breakdown voltage    ProcessbvV0      o     s����� 1.0e-3$Current at reverse breakdown voltage    ProcessibvA0      p     s�����  Ohmic conductance    ProcesscondMho     r        D��     m���                Ariald     h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  COpAnal                         
                        ����            ���               ��  TSignal                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                      v(iv_vl)       ����                  n�	                     	i(va_ix1)       ����                  n�
                     i(va_il)       ����                  n�                      	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CDCsweep       
 3456789:;<               
                       ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                       v(iv_vl)       ����                  n�	                      	i(va_ix1)       ����                  n�
                      i(va_il)       ����                  n�                       	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACsweep        MNOPQRST               
                       ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                      v(iv_vl)       ����                  n�	                     	i(va_ix1)       ����                  n�
                     i(va_il)       ����                  n�                      	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  �� 
 CTranSweep       klmnopqr               
                       ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                       v(iv_vl)       ����                  n�	                      	i(va_ix1)       ����                  n�
                      i(va_il)       ����                  n�                       	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACdisto        fghij               
                           ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                       v(iv_vl)       ����                  n�	                      	i(va_ix1)       ����                  n�
                      i(va_il)       ����                  n�                       	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��        #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
                          ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                       v(iv_vl)       ����                  n�	                      	i(va_ix1)       ����                  n�
                      i(va_il)       ����                  n�                       	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��        #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
                           ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                       v(iv_vl)       ����                  n�	                      	i(va_ix1)       ����                  n�
                      i(va_il)       ����                  n�                       	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��        #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
                           ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                       v(iv_vl)       ����                  n�	                      	i(va_ix1)       ����                  n�
                      i(va_il)       ����                  n�                       	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��        #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
                           ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                       v(iv_vl)       ����                  n�	                      	i(va_ix1)       ����                  n�
                      i(va_il)       ����                  n�                       	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��        #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
         2             	    ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                      v(iv_vl)       ����                  n�	                     	i(va_ix1)       ����                  n�
                     i(va_il)       ����                  n�                      	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACnoise        UVWXYZ[\               
                    
    ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                      v(iv_vl)       ����                  n�	                     	i(va_ix1)       ����                  n�
                     i(va_il)       ����                  n�                      	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  �         #�  ����        ��������#�  ����       ��������#�  ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������              
                        ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                      v(iv_vl)       ����                  n�	                     	i(va_ix1)       ����                  n�
                     i(va_il)       ����                  n�                      	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CFourier        stuv               
         ��                   ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                      v(iv_vl)       ����                  n�	                     	i(va_ix1)       ����                  n�
                     i(va_il)       ����                  n�                      	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACpz        	 ]^_`abcde               
                       ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                      v(iv_vl)       ����                  n�	                     	i(va_ix1)       ����                  n�
                     i(va_il)       ����                  n�                      	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CDCtf         =>?@A               
                       ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                      v(iv_vl)       ����                  n�	                     	i(va_ix1)       ����                  n�
                     i(va_il)       ����                  n�                      	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CDCsens         BCDEFGHIJKL               
                       ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                       v(iv_vl)       ����                  n�	                      	i(va_ix1)       ����                  n�
                      i(va_il)       ����                  n�                       	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j                  ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                      v(iv_vl)       ����                  n�	                     	i(va_ix1)       ����                  n�
                     i(va_il)       ����                  n�                      	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CShow         w              
                       ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                      v(iv_vl)       ����                  n�	                     	i(va_ix1)       ����                  n�
                     i(va_il)       ����                  n�                      	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CShowmod         x              
                       ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                      v(iv_vl)       ����                  n�	                     	i(va_ix1)       ����                  n�
                     i(va_il)       ����                  n�                      	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  �� 
 CLinearize        #�  ����        ��������               
                       ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                      v(iv_vl)       ����                  n�	                     	i(va_ix1)       ����                  n�
                     i(va_il)       ����                  n�                      	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CParamTranSweep        yz{|}~������               
                       ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                      v(iv_vl)       ����                  n�	                     	i(va_ix1)       ����                  n�
                     i(va_il)       ����                  n�                      	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  |              ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                       v(iv_vl)       ����                  n�	                      	i(va_ix1)       ����                  n�
                      i(va_il)       ����                  n�                       	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CParamACSweep        ����������                
                       ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                      v(iv_vl)       ����                  n�	                     	i(va_ix1)       ����                  n�
                     i(va_il)       ����                  n�                      	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CMonteCarlo_op        ����������������������������               
                              ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                      v(iv_vl)       ����                  n�	                     	i(va_ix1)       ����                  n�
                     i(va_il)       ����                  n�                      	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CMonteCarlo_dc        ����������������������������               
                       ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                       v(iv_vl)       ����                  n�	                      	i(va_ix1)       ����                  n�
                      i(va_il)       ����                  n�                       	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CMonteCarlo_ac        ����������������������������               
                       ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                      v(iv_vl)       ����                  n�	                     	i(va_ix1)       ����                  n�
                     i(va_il)       ����                  n�                      	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CMonteCarlo_tran        ����������������������������               
                       ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                       v(iv_vl)       ����                  n�	                      	i(va_ix1)       ����                  n�
                      i(va_il)       ����                  n�                       	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACsens        	
               
                              ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                       v(iv_vl)       ����                  n�	                      	i(va_ix1)       ����                  n�
                      i(va_il)       ����                  n�                       	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CNetworkAnalysis                       
                       ����            P               n�                        v(ctrl)       ����                  n�                       v(13)       ����                  n�                       v(3)       ����                  n�                       v(4)       ����                  n�                       v(5)       ����                  n�                       v(9)       ����                  n�                       v(11)       ����                  n�                       i(v1)       ����                  n�                       v(iv_vl)       ����                  n�	                      	i(va_ix1)       ����                  n�
                      i(va_il)       ����                  n�                       	v(iv_vx1)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j                  ����            P                 >           ��   CDigSimResTemplate                ���       ����  ����:�0�yU>20.00n���   ����                       Arial����                       Arial����                       Arial  �   �  �                                ����  ���� ������       ����  ���� ������                 �               ����  �����       200������         0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial      �       �         �     �   �  �  Circuit1                  ����  ��    ��������                                                                                                                                                                           g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     ��   CPackageAliasSuperPCBStandardDIODE3      �Eagle	DIODE.LBRDO41-7   AC  �Orcad 	DAX2/DO41      �	Ultiboard	L7DIO.l55DIO_DO41              A                                                            g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     �SuperPCBStandardDIODE3      �Eagle	DIODE.LBRDO41-7   AC  �Orcad 	DAX2/DO41      �	Ultiboard	L7DIO.l55DIO_DO41              A                                                g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     �SuperPCBStandardDIODE3      �Eagle	DIODE.LBRDO41-7   AC  �Orcad 	DAX2/DO41      �	Ultiboard	L7DIO.l55DIO_DO41              A      g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     �SuperPCBStandardDIODE3      �Eagle	DIODE.LBRDO41-7   AC  �Orcad 	DAX2/DO41      �	Ultiboard	L7DIO.l55DIO_DO41              A                                                          �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D  �                . C�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                      �  �                �         �  @                  ���                                                  �  @  �     <   �  <     ��                                                        �     |   �  |     ��                                                        �     �   �  �     ��                                                        �     �   �  �     ��                                                        � �      �  4     ��                                                      �      �  4   �      �  4   [title]                                       � �   D   �  t     ��                                                      �   D   �  t   �   D   �  t   [description]                                       � `   �   h  �     ��                                                      `   �   h  �   `   �   h  �   [id]                                       � �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       �      �   8    ��        	                                                   �   8       �   8  Date :       �    H
  �                  � �     �  4   	 ��        
                                              �     �  4  �     �  4  [date]                                       �       t   8    
 ��                                                            t   8         t   8   Title :       �     
  �                  �    L   �   x     ��                                                         L   �   x      L   �   x   Description :       �  �  �  �                  �    �   �   �     ��                                                         �   �   �      �   �   �   ID :       �  �  �	  P                  �    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �  \  8                     012345678:;<=>          9     	title box    Analog Misc      �?    9 
 l�     #�  ����        ��������#�  ����       ��������#�  ����       ��������#�  ����       ��������#�  ����       ��������        9                                      ����q��� ����     s�            title                s�            description               s�            id               s�            designer               s�            date                           ����            `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                                                                                            2         �  �              � � �                   ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                          �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   
cgs 76         47 80moh5.6 ���� � mvrd nmodel            
 n�                      TIME� # ) time                      n�                        i(v1)� < � i(v1)    TIME                 n�                        v(3)      v(3)    TIME                 n�                      	i(va_ix1)�   � 	i(va_ix1)    TIME                 n�    (v(7)-v(3))                   v(IV_VL)� �   v(IV_VL)    TIME                 n�                      i(va_il)  � � i(va_il)    TIME                 n�    v(5)                   	v(IV_Vx1)� �   	v(IV_Vx1)    TIME                 n�    v(iv_vx1)*i(va_ix1)                    Pin� # )  ����TIME                 n�                       v(ctrl)      v(ctrl)    TIME                 n�                        v(5)      v(5)    TIME                           2         �  �           Time  � � �                   ����                       Arial����                       Arial                              ����  ������}���?1.539715e-002��k-	      ����  �����ZE8�Zs?4.725051e-003��M��      ����  ����]�P�N@5.576897e+000������      ����  �������9���-1.971735e+000������                                                                         �                      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �  �                                                                                                                                                                                                                                                                                                                                                                                                                                  �
  �
                                                                      �  �                                                                      �  �                                              1m  0                            100   100                                                             1m  0                            100   100                                1m  0                            100   100                                1m  0                            100   100                                                 
                 1m  0                            100   100                            ��   CPartPackage     ��   CPackageg   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     *+,-   W��/� Y�g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     &'()   W�     Y�g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     "#$%   W���� Y�g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �      !      ��   CMiniPartPin    ����V+V+     PWR+V+g      a�   ����V-V-     PWR-V-h     voltage_sourcevoltage_source                          a�    ����C+C+     PASC+�      a�   ����C-C-     PASC-�     capacitor_genericcapacitor_generic                          a�    ����11     PAS1�      a�   ����22     PAS2�     BatteryBattery                          a�    ����R+R+     PASR+      a�   ����R-R-     PASR-     RR                          a�    ����GndGnd     GNDGnd}      GndGnd                  a�    ����M+M+     PASM+i      a�   ����M-M-     PASM-j     	voltmeter	voltmeter                          a�    ����M+M+     PASM+2      a�   ����M-M-     PASM-3     Ammeter2Ammeter2                          a�    ����GndGnd     GNDGnd}      GndGnd                  a�    ����GndGnd     GNDGnd}      GndGnd                  a�    ����MM       ��������MarkerMarker                  a�    ����GndGnd     GNDGnd}      GndGnd                  a�    ����MM       ��������MarkerMarker                  a�    ����MM       ��������MarkerMarker               _ a�    ����D+D+     PASA       a�   ����D-D-     PASK       !  ��   CPackagePin 1 D+PAS  AAw� 2 D-PAS  AKDiodeDiode	Fairchild      1n4007 D1n4007D4            diode-21n40071n4007                          a�    ����GndGnd     GNDGnd}      GndGnd                  a�    ����11     PAS1S      a�   ����22     PAS2T     a�   ����33     PAS3U     a�   ����44     PAS4V     vcswitchvcswitch                                          a�    ����GndGnd     GNDGnd}      GndGnd                  a�    ����MM       ��������MarkerMarker               ] a�    ����D+D+     PASA       a�   ����D-D-     PASK       �  w� 1 D+PAS  AAw� 2 D-PAS  AKDiodeDiode	Fairchild      1n4007 D1n4007D3            diode-21n40071n4007                          a�    ����L+L+     PASL+K      a�   ����L-L-     PASL-L     InductorInductor                          a�    ����M+M+     PASM+0      a�   ����M-M-     PASM-1     AmmeterAmmeter                          a�    ����M+M+     PASM+k      a�   ����M-M-     PASM-l     
Voltmeter2
Voltmeter2                       [ a�    ����D+D+     PASA       a�   ����D-D-     PASK       Q  w� 1 D+PAS  AAw� 2 D-PAS  AKDiodeDiode	Fairchild      1n4007 D1n4007D2            diode-21n40071n4007                       X a�    ����D+D+     PASA       a�   ����D-D-     PASK       W  w� 1 D+PAS  AAw� 2 D-PAS  AKDiodeDiode	Fairchild      1n4007 D1n4007D1            diode-21n40071n4007                          a�    ����11     PAS1S      a�   ����22     PAS2T     a�   ����33     PAS3U     a�   ����44     PAS4V     vcswitchvcswitch                                          a�    ����11     PAS1S      a�   ����22     PAS2T     a�   ����33     PAS3U     a�   ����44     PAS4V     vcswitchvcswitch                                          a�    ����11     PAS1S      a�   ����22     PAS2T     a�   ����33     PAS3U     a�   ����44     PAS4V     vcswitchvcswitch                                                                                                                                                                                                    
m1     8 8 mm l=100u w                        used                            ��    �Z�P��,�                        ��                                                                                                            (f    x=f � �'f                           �(f                            ,�e    �f � ��e                           ��e                                     �  � ���� �                         .I                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       h�    ���������                        ��                            @R    �`R``R�_Rx_R                        pbR                                                                                                            �$�    h&��&��&� '�                        H)�                            MJ         W X Y [   Z                          DIN                            sist      resistor DIN                                                       ��S    ��S0�S��S��S                        �S                            ��    ��������P��                        ��                            �V�    (W�`W��W��W�                        �Y�                            Їl    `�l(�l`-j �W                         �W                            t�@
    L �k��
>ENDDATA
                        
JV1                            p�<        ��<x�                           �                                                                                                                                                                                            �2�    �Q�R�XR��R�                        T�    2 2 2 2 d                                                                                                         