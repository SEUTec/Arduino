    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz    ��  CPart    �����   �  �  �����   �  �              voltage_source��  CIntPin    ��  CWire    �        �
   /   �   �      /   �   �                  Marker ��  CExtPin    ��  CVertex
   �      ��  CSegment;    �G   �  `                 �:    �Q   �      �/    �"   �  `                           
        `      M     �  �          Ctrl     ��   CPin                   ��                                                           `   M��  TLine     P       `     ��    ��                                                ��  TPolygon     ����    ����   ��                                                         ��  TPoint    0        �   @        �    P        �0   @            ��  
 TTextField    �����        ��                                                          �����         �����      	[refname]       �  �  8  g        �   ,                Marker     Miscellaneous      �?    +   ��   CMarkerBehavior     ��  CValue ����    �i��       �������� M ��  	 TModelPin ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      "   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               & Analog MiscV   Generic   CtrlCtrl          ����               Ctrl  v(Ctrl)  N ��   CPartPin    ����MM       A H� ����RootmarkerGeneric              Ctrl  �      �       �   �  �      �   �  �              vcswitch�    �    �    ,   �       _   �         _   �                 capacitor_generic- �   �    / �   0   �       S   �  ,      S   �  ,              Ammeter�    �    �   4   �       �   �        �   �                Inductor�    �    �    8    �       �   �  �       �   �  �               R9 �   ,   : 3 	�    �    
  �	   �8   = �   @  �	   >                        �  �   R+  	�   �   �  �	   �9   �P   �  �	   B �   �5   �  @   �    E �8    
  @   F            D �   �O   �  �   �5   I �   @  �   J             �   �>   �  �   L         I     H     E         C     �   �F   �  �   N        C         A                  �   R-   �   	         R     �                    ��                                                       �   @   R+�                   ��                                                          @   R-�    @   $   0     ��    ��)                                                � 0   P   $   0     ��                                                        � 0   P   <   0     ��    ��)                                                � H   P   <   0     ��    p�Z                                                � H   P   T   0     ��                                                       � `   P   h   @     ��    D�Z                                                � �   @   h   @     ��    ��d                                                � `   P   T   0    	 ��    |�f	                                                �    @       @    
 ��    <�b
                                                �     `   �   �     ��                                                           `   �   �       `   �   �   [resistance]       �   
  `	  �
      `   �   �   �         t   $     ��                                                               t   $           t   $   	[refname]       �   	  �  �	          t   $    P Q R S T U V W X Y Z [ \    resistor    resistor DINMiscellaneous      �?       ��  CResistorBehavior     #� �������(\��?0.58      ��������#� ���� 27     ��������#� ����       ��������#� ����       �������� R+R- ��   CBehPin     R+        ����R+����                        ��c�    R-      ����R-����                        �� resistor                d e Passive   Generic   RR          ����    R '�    ����R+R+      PASAR+    ����'�   ����R-R-      PASAR-    ����Passivedefault resistor, 1KGeneric              5 7  d c�     L+        ����L+����                        �� 5   6 5 5 	�    ?        �   L+K  	�   �      �	   �6   k �.   �  �	   l                      �  �   L-L   @   	          L1     �                    ��                                                           @   L+�                   ��                                                      �   @   L-��   TArc h   ,   �   T    
                                                           h   ,   �   T   h   ,   �   T   �   @   h   @           p� P   ,   h   T    	                                                           P   ,   h   T   P   ,   h   T   h   @   P   @           p� 8   ,   P   T                                                               8   ,   P   T   8   ,   P   T   P   @   8   @           p�     ,   8   T                                                                   ,   8   T       ,   8   T   8   @       @           � $   P      X     ��    ��                                                �    H   $   P     ��     �                                                  �     P   $   P     ��    ��                                                �     @       @     ��    p�H	                                                � �   @   �   @     ��       
                                                �     \   �   |     ��                                                           \   �   |       \   �   |   [Inductance]       @  
  @  �
      \   �   |   �         �   $     ��                                                               �   $           �   $   	[refname]       @   	  �  �	          �   $    n o y   x   w   v   u z {   t   s   r   q      Inductor     Miscellaneous      �?    
   ��  CInductorBehavior     #� ��� �������?100m      ��������#� ���� x     �������� L+L- h c�    L-      ����L-����                        �� Inductor  
              h � Passive   Generic   L1L1          ����  L '�    ����L+L+      PASAL+������'�   ����L-L-      PASAL-�D� ����PassiveInductorGeneric              11 3  � c�     M+        ����M+����                        �� 11   2 11 1 	�    m        �   M+0  	�   �   �  �	   �3   � �I   @  �	   � �   � �)   @  �   �            �   �A   @  @   �-   �%      @   �         �     � �%   �C   @  �   �(   �-   �  �   �        �     �+   �9   @  �   �         �     �     �         �                      �  �   M-1   �   	          VA_IL    	 �                   ��                                                           @   M+�                   ��                                                      �   @   M-� �   @   �   @     ��    ��                                                �     @       @     ��                                                        � 4   X   `   X     ��    ��                                                �� 
 TRectangle        �   d                   ����                                                �   d   � ����������������  ��          @ @                                           �d   X    IX1.�X   P        �X   `    0000@ @ � $   $   �   L     ��                                                      $   $   �   L   $   $   �   L   [value]                       $   $   �   L   �     �����        ��                                                           �����          �����      	[refname]       @  �  X  r	      �����       �   � � �   �   � � �   � 	     Ammeter    Ammeter_smallMiscellaneous      �?       ��   CAmmeterBehavior     #� ����    �i��       �������� M+M- � c�    M-      ����M-����                        ��AmmeterAmmeter   �            � � Analog Meters   Generic   VA_ILVA_IL          ����  VAm '�    ����M+M+      PASAM+XQ� ����'�   ����M-M-      PASAM-�R� ����Analog MetersAmmeterGeneric              13 �   0   �       �   �  �      �   �  �              vcswitch�    �     �    �     �           �   �           �   �               Gnd� 	�    �+   `  `   �<   �   `  `	   �         �     �*   �J      `   �4   �      @   �         �     �      �     �$   � �?   �  `   �)   �L   �  �   �          �     � �   � �;   @  `   �&   �M   @  @   �'   �<   @  �   �      �     �          �     �                               `       Gnd}      `          gnd1     �                    ��                                                               Gnd�                   ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��    p�Z         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         � � � �   �      Ground    
Ground DINMiscellaneous      �?       ��   CGroundBehavior       Gnd c�     Gnd        ����Gnd����                        ��gndgnd                 � Analog Meters   Generic   gnd1gnd1          ����  gnd '�    ����GndGnd      GNDAGnd �)����SourcesGroundGeneric              0 �   �    �           �   �          �   �              Battery�    �    � �    �    �       _   @  �      _   @  �              Ammeter2� �   �    � �    �    �       _   �  �      _   �  �              
Voltmeter2� �   �    � 0 	�    �(      �   �,   �@      �    � �   � �H   `  �    �2   � �   `  �   �            � �"   � �D   �  �    �.   � �#   �  `   �            � �!   � �:   @  �    � �#   � �B   @  `   �                                        �                `   `   M+k  	�   �   `   �  M-l   �   `          IV_Vx1    
 �                    ��                                                               M+�                   ��                                                          �   M-�     �       �     ��    ��                                                �             <     ��    
NVA                                                �    $      4     ��    ��                                                �    ,      ,     ��    p�H                                                �    �      �     ��               	FIXED_ROT                                        ��     <   �   �                  ����                                             <   �   �   �    D   �   x     ��                                                         D   �   x      D   �   x   [value]                          D   �   x   � 8      �   0    	 ��        	                                               8      �   0   8      �   0   	[refname]       h  �  �    8      �   0    � � � � � � �     �       �   � 
     Voltemeter-Vert    Voltemeter-Vert_smallMiscellaneous      �?       ��   CVoltmeterBehavior     #� ����    �i��       �������� M+M- c�     M+        ����M+����                        ��c�    M-      ����M-����                        ��	voltmeter	voltmeter   k            � � Analog Meters   Generic   IV_Vx1IV_Vx1          ����  IVm '�    ����M+M+      PASAM+   ����'�   ����M-M-      PASAM-�tc����Analog MetersVoltmeter-verticalGeneric              9 �   �   * 9 �   �   �       �   �         �   �                 1n4007�    0    � 13 � 	�    �        @  D+   	�   �          D-    @  @         D1     �                   ��                                                           �   D+�                   ��                                                          `   D-� �����       �      ��    ���                                                 �     �       �     ��                                                        � �����       �     ��    ���                                                 �     �       �     ��    (�K                                                � �����       �     ��                                                       �     �      �     ��    ��K                                                �     �       `     ��    ��K                                                � d   �   $  �    	 ��        	                                               0   `   �   �   0   `   �   �   	[devname]        �������������������������      � 0   �   �   �    
 ��        
                                               0   �   �   �   0   �   �   �   	[refname]       �  �  P  �  ����   �   <    � �                � �  �
  diode     Miscellaneous      �?       ��  CDiodeBehavior     #� ����        ��������#� ���� 27     ��������#� ����       ��������#� ����       �������� D+D- c�     D+        ����D+����                        ��c�    D-      ����D-����                        ��d1n4007d1n4007    �          Diode   Generic   D1D1                D '�    ����D+D+      PASAA�נ ����'�   ����D-D-      PASAK(٠ ����DiodeDiode	FairchildDO-41             9  c�    M-      ����M-����                        ��c�    2      ����2����                        ���  9  � 9 	�    �   `  `   �7   �   `  �                          `   �  M+2  	�   �   `   `   M-3      �         VA_Ix1    	 �                    ��                                                           �   M+�                   ��                                                              M-�     �       �     ��                                                        �     <             ��                                                        �� @   <   �����                  ����                                         ����<   @   �   � ����x   ����L     ��                                                        �  ������� �������  ��          @ @                                           �����H    ��b�����T    
>DA�����T    uT@ @ � ����D   <   |     ��                                                      ����D   <   |   ����D   <   |   [value]                          D   �   |   � ��������O        ��                                                       ��������O      ��������O      	[refname]       �  _  �  �     �����      
 "  #	   Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       ��     #� ����    �i��       �������� M+M- c�     M+        ����M+����                        ��AmmeterAmmeter   V            &Analog Meters   Generic   VA_Ix1VA_Ix1          ����  VAm '�    ����M+M+      PASAM+ '����'�   ����M-M-      PASAM-�� ����Analog MetersAmmeter-verticalGeneric              4  c�     1       ����1����                        ��& 4   � 4 � 	�       `       1�  	�   �   `   �  2�      �          XSource     �                    ��                                                               1�                   ��                                                          �   2�             $     ��    ��)                                                �     \       �     ��                                                        �    8   0   8    	 ��    ��)                                                �     H   @   H     ��    p�Z                                                �     $   @   $     ��                                                       �    \   0   \     ��    D�Z                                                �               ���                                                      �               ���   �Z	                                                � `          $    
 ��        
                                               `          $   `          $   	[devname]        ����������������`          $   � `   $      H     ��                                                       `   $      H   `   $      H   	[refname]          L  �  �  `   $      H    ,-./2345    67    1  0     Battery     Miscellaneous      �?    9 
 ��  CParamSubBehavior     #� ����      (@12      �������� 12 )c�    2      ����2����                        ��BatteryBattery
 9 i             );Sources   Generic   XSourceXSource          ������   CParamSubModelType��    BATTERY2.SUBCKT Xbattery 1 2
V1 1 2 DC {voltage}
.ENDS
   ��  	 CParmDefn    1battery voltage   ParamSubvoltageV                X '�    ����11      PASA1    ����'�   ����22      PASA2 � ����SourcesBatteryGeneric              0 � �    �     �       �   �         �   �                 1n4007B�   ,   C3 	�    �        @  D+   	�   O          D-    �  �         D2     �                   ��                                                           �   D+�                   ��                                                          `   D-� �����       �      ��    ���                                                 �     �       �     ��                                                        � �����       �     ��    ���                                                 �     �       �     ��                                                       � �����       �     ��    ��K                                                �     �      �     ��    ��K                                                �     �       `     ��                                                        � d   �   $  �    	 ��        	                                               0   `   �   �   0   `   �   �   	[devname]        �������������������������      � 0   �   �   �    
 ��        
                                               0   �   �   �   0   �   �   �   	[refname]         \  �  �  ����   �   <    IJKLMNO    PQ          GH �
  diode     Miscellaneous      �?       �     #� ����  F      ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     �������� D+D- c�     D+        ����D+����                        ��c�    D-      ����D-����                        ��d1n4007d1n4007    @          WXDiode   Generic   D2D2                D '�    ����D+D+      PASAAb����'�   ����D-D-      PASAK�b����DiodeDiode	FairchildDO-41             0 � �    �     �           �   �           �   �               Gnd[	�    �   �  �                     `       Gnd}   �  �          gnd4     �                    ��                                                               Gnd�                   ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��    D�H         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��    x�W         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��    X��         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         _`ac  b     Ground    
Ground DINMiscellaneous      �?       ŀ       Gnd c�     Gnd        ����Gnd����                        ��gndgnd                 eAnalog Meters   Generic   gnd4gnd4          ����  gnd '�    ����GndGnd      GNDAGndP�e����SourcesGroundGeneric              0 �   �     0 �    �     �           �   �           �   �               Gndh	�    �   �  �                    `       Gnd}   `  �          gnd5     �                    ��                                                               Gnd�                   ��    p�H         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��    D�H         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         lmnp  o     Ground    
Ground DINMiscellaneous      �?       ŀ       Gnd c�     Gnd        ����Gnd����                        ��gndgnd                 rAnalog Meters   Generic   gnd5gnd5          ����  gnd '�    ����GndGnd      GNDAGnd�9b����SourcesGroundGeneric              0 �   �    * 0 �    �     �           �   �           �   �               Gndu	�    �      @                    `       Gnd}   �  @          gnd6     �                    ��                                                               Gnd�                   ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��       0         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��       �         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         yz{}  |     Ground    
Ground DINMiscellaneous      �?       ŀ       Gnd c�     Gnd        ����Gnd����                        ��gndgnd                 Analog Meters   Generic   gnd6gnd6          ����  gnd '�    ����GndGnd      GNDAGnd Bb����SourcesGroundGeneric              0 �   �    � 0 �    �     �           �   �           �   �               Gnd�	�    �K   �  @                    `       Gnd}      @          gnd7     �                    ��                                                               Gnd�                   ��     �          AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��    @�Y         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��    X�Y         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��    X�Z         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         ����  �     Ground    
Ground DINMiscellaneous      �?       ŀ       Gnd c�     Gnd        ����Gnd����                        ��gndgnd                 �Analog Meters   Generic   gnd7gnd7          ����  gnd '�    ����GndGnd      GNDAGnd�db����SourcesGroundGeneric              0 �   �    �   �����   �  �  �����   �  �              voltage_source�    �    �    �   �   /   �   �      /   �   �                  Marker�	�    �      `   �1   ��E   �  `   ��   ��N   �  �   �                    �0   ��!      �   �                      `      Mhz� �  @          Ctrl2     �                   ��                                                           `   M�     P       `     ��                                                        �     ����    ����   ��                                                         �    0        �   @        �    P        �0   @            �    �����        ��                                                          �����         �����      	[refname]       �  1  �  �        �   ,    �  ���     Marker     Miscellaneous      �?    +   !�     #� ����    �i��       �������� M %� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     ��  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               �Analog MiscV   Generic   Ctrl2Ctrl2          ����               Ctrl2  v(Ctrl2)  N '�    ����MM       A ��������RootmarkerGeneric              Ctrl2 ��   �  � Ctrl2  �c�    3      ����3����                        ��c�     V+        ����V+����                        �� Ctrl2   �Ctrl2 �	�    �          V+g  	�   �      �  V-h   �  �         V2     �                   ��                                                           `   V+�                   ��                                                          �   V-��  TEllipse     �   �����                   ����                                         �����       �   �����       �   �    �   �����     ��    V                                                �     �       �     ��    `                                                   �     �       �     ��     �                                                 �     \       �     ��                                                        � �����   
   �    
 ��                	FIXED_ROT                                        � \   `   \   `     ��                                                      \   `   \   `   \   `   \   `           �  �  �  �                � 0   �   �   �     ��        	                                               0   �   �   �   0   �   �   �   [dc]         P  H  �          p   @   � 0   \   �   �    	 ��        
                                               0   \   �   �   0   \   �   �   	[refname]         �  �  J      ����t       �  ��������      �    � �  Voltage Source    Voltage Source DINRoot      �?       ��  CVSourceBehavior     #� ����        0      ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       �������� V+V- �c�    V-      ����V-����                        ��volt_sourcevolt_source   +0            ��Sources   Generic   V2V2          ����       #�0            0      ��������#�0����      @5     ��������#�0            0     ��������#�0'  ���ư>1u     ��������#�0'  ���ư>1u     ��������#�0 -1����Mb`?2m     ��������#�0 '�~j�t��?12m     ��������    #�0            0      ��������#�0����      �?1.5     ��������#�0����      I@50     ��������#�0            0     ��������#�0            0     ��������    #�0            0      ��������#�0����      �?1     ��������#�0����      �?1     ��������#�0            0     ��������#�0����      �?1     ��������    #�0            0      ��������#�0����      �?1     ��������#�0            0     ��������#�0 N  �����>2u     ��������#�0'  ���ư>1u     ��������#�0'  ���ư>1u     ��������    #�  ���� 0 0      ��������                0      �������� ����       �������� ����       �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������               V '�    ����V+V+      PWR+AV+p�b����'�   ����V-V-      PWR-AV- 1b����Sources Generic              0  c�    V-      ����V-����                        ��;� erc�    4      ����4����                        ��� W�c�     1       ����1����                        ��c�    4      ����4����                        ���  0    � 0 � ��	�    �        �  1S  	�   �          2T  	�   �  �      3U  	�   x  �   �  4V   @  �         X2     �                    ��                                                           �   1�                   ��                                                          `   2�                   ��                                                      @   `   3�                   ��                                                      @   �   4� @   �   @   �     ��    ���                                                 � @   `   @   �     ��    |-S                                                � @   �   @   �    
 ���   ���                                                 � H   �   8   �    	 ���   (�K                                                ��    �   �����                  ����                                         �����      �   �����      �   �� P   �   0   �               	   ����                                         0   �   P   �   �     `       �     ��       
                                                �    �       �     ��    ��K                                                �     �       �     ��                                                       � 8   �   H   �     ��  � ԎK        	FIXED_ROT                                        � ,   �      �     ��                                                        � `   �   �   �     ��                                                       `   �   �   �   `   �   �   �   	[refname]       `  \  �  �      (   t   L   � `   `   �   �     ��                                                       `   `   �   �   `   `   �   �   	[devname]        ����������������       �   (    �������      ��  �������    � �  vcswitch     Miscellaneous      �?   9 
 8�    #� ����      �?1      ��������#� ������������-1.3     ��������#� ����      �?0.5     ��������#� ����    ��.A1meg     �������� 1234 �c�    2      ����2����                        ����X5_vcswitchX5_vcswitch
 9               � ��Switches   Generic   X2X2          ����<���voltage controlled switch   VCSW{.subckt vcsw 1 2 3 4
S 1 2 3 4 switch
.model switch sw (vt={(Von+Voff)/2} vh={(Von-Voff)/2} ron={Ron} roff={Roff})
.ends   >�    1turnon voltage   ParamSubVon               >�    1turnoff voltage   ParamSubVoffV             >�    0on resistance   ParamSubRonOhm             >�    0off resistance   ParamSubRoffOhm               X '�    ����11      PASA1G4  ����'�   ����22      PASA2    ����'�   ����33      PASA3� b����'�   ����44      PASA4�އ ����Switches Generic              13 �   0   �       �   �  �      �   �  �              	voltmeter�    ,    3 
	�    K           M+i  	�   �   �     M-j   @  �          IV_VL    
 �                   ��                                                           `   M+�                   ��                                                      �   `   M-�     `       `     ��    ��                                                � �   `   �   `     ��                                                        �    L      \     ��    ��                                                �     T      T     ��    p�H                                                � �   X   �   X     ��               	FIXED_ROT                                        ��     <   �   �                   ����                                             <   �   �   � (   D   �   x     ��                                                      (   D   �   x   (   D   �   x   [value]                       (   D   �   x   �        �   0    	 ��        	                                                      �   0          �   0   	[refname]       �  �  �  Z         �   0              
     	voltmeter    voltmeter_smallMiscellaneous      �?       �     #� ����    �i��       �������� M+M- c�     M+        ����M+����                        ��c�    M-      ����M-����                        ��	voltmeter	voltmeter   _            Analog Meters   Generic   IV_VLIV_VL          ����  IVm '�    ����M+M+      PASAM+c����'�   ����M-M-      PASAM-X#c����Analog Meters Generic              13 �  c�    C-      ����C-����                        ���   13   . 13 	�    �   �  �   C-�  	�   G        �   C+�    
  �          C1     �                   ��                                                       �   @   C-�                   ��                                                          @   C+�     @   @   @      ��    ���                                                 � @       @   `     ��    �b�                                                � `       `   `     ��    ���                                                 � `   @   �   @     ��    (�K                                                �     `   �   �     ��                                                           `   �   �       `   �   �   [capacitance]        
  �  �
  ,	      `   �   �   �         �   $     ��                                                               �   $           �   $   	[refname]        
  �  �
            �   $    $%&'(    )      "#     	Capacitor     Miscellaneous      �?       ��  CCapacitorBehavior     #� '  �dy���=20p      ��������#� ���� x     ��������#� ����       ��������#� ����       �������� C+C- c�     C+        ����C+����                        �� 	capacitor                0Passive   Generic   C1C1          ����  C '�    ����C+C+      PASAC+�-c����'�   ����C-C-      PASAC-8/c����Passive Generic              3 ; D+  0e c�     1       ����1����                        ��X 3   * 3 � ) t	�    M    �   �  1S  	�   �   �      2T  	�             3U  	�   k      �  4V   �  @        X1     �                    ��                                                       @   �   1�                   ��                                                      @   `   2�                   ��                                                          `   3�                   ��                                                          �   4�     �       �     ��                                                        �     `       �     ��                                                        �     �       �    
 ���                                                       � �����      �    	 ���                                                       �� D   �   <   �                  ����                                         <   �   D   �   <   �   D   �   ��    �   �����               	   ����                                         �����      �   � @   `   @   �     ��        
                                                � 0   �   @   �     ��                                                        � @   �   @   �     ��                                                        �    �   �����     ��  �             	FIXED_ROT                                        �    �   4   �     ��                                                        � `   �   �   �     ��                                                       `   �   �   �   `   �   �   �   	[refname]       �  �  P  �      (   t   L   �     �  <    ��                                                       `   `   �   �   `   `   �   �   	[devname]        ����������������       �   (    89:;ABD      =E  F?GHC<>    @ �  vcswitch     Miscellaneous      �?   9 
 8�    #� ����      �?1      ��������#� ����      �?1     ��������#� ����      �?0.5     ��������#� ����    ��.A1meg     �������� 1234 3c�    3      ����3����                        ���X6_vcswitchX6_vcswitch
 9               3N�Switches   Generic   X1X1          ����<���voltage controlled switch   VCSW{.subckt vcsw 1 2 3 4
S 1 2 3 4 switch
.model switch sw (vt={(Von+Voff)/2} vh={(Von-Voff)/2} ron={Ron} roff={Roff})
.ends   >�    1turnon voltage   ParamSubVon               >�    1turnoff voltage   ParamSubVoffV             >�    0on resistance   ParamSubRonOhm             >�    0off resistance   ParamSubRoffOhm               X '�    ����11      PASA1p�b����'�   ����22      PASA2(yc����'�   ����33      PASA3�އ ����'�   ����44      PASA4��b����Switches Generic              Ctrl  c�     V+        ����V+����                        ��& N Ctrl    Ctrl g	�               V+g  	�   ^      �  V-h   �  @         V1     �                   ��                                                           `   V+�                   ��                                                          �   V-��     �   �����                   ����                                         �����       �   �����       �   �    �   �����     ��    ��)                                                �     �       �     ��    ��`                                                �     �       �     ��    ��)                                                �     \       �     ��    p�Z                                                � �����   
   �    
 ��               	FIXED_ROT                                        � \   `   \   `     ��                                                      \   `   \   `   \   `   \   `           �  `  �  `                � 0   �   �   �     ��        	                                               0   �   �   �   0   �   �   �   [dc]       p  �  �  |          p   @   � 0   \   �   �    	 ��        
                                               0   \   �   �   0   \   �   �   	[refname]       p  T  �  �      ����t       ]  ^_a\`cde      b    [ �  Voltage Source    Voltage Source DINRoot      �?       ��     #� ����        0      ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       �������� V+V- X�volt_sourcevolt_source   +0            X�Sources   Generic   V1V1          ����       #�0            0      ��������#�0����      @5     ��������#�0            0     ��������#�0'  ���ư>1u     ��������#�0'  ���ư>1u     ��������#�0 -1����Mb`?2m     ��������#�0 '�~j�t��?12m     ��������    #�0            0      ��������#�0����      �?1.5     ��������#�0����      I@50     ��������#�0            0     ��������#�0            0     ��������    #�0            0      ��������#�0����      �?1     ��������#�0����      �?1     ��������#�0            0     ��������#�0����      �?1     ��������    #�0            0      ��������#�0����      �?1     ��������#�0            0     ��������#�0 N  �����>2u     ��������#�0'  ���ư>1u     ��������#�0'  ���ư>1u     ��������    #�  ���� 0 0      ��������                0      �������� ����       �������� ����       �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������               V '�    ����V+V+      PWR+AV+NDDA����'�   ����V-V-      PWR-AV- � ����Sources Generic              . � : � �        \        i* v�      6 2 � � C�� �	 	 	 �  �0 , � 8 � 4 = & =                                     �  �     N H   � D L   � � F � � � � � � � � � � � � � �  ��� � � J l > B   � R 3 R   � ^               x  k  A =   k ?       K �   �   � �  � �   �     � �   �   � m             E     G � � � �   M � � � � � � �O  � � � �� � �I C     ��  CLetter    �Los dos interruptores se ponen en ON al mismo tiempo.
X2 se pone en OFF, deja de fluir corriente desde la fuente.
Entonces la corriente retorna a la fuente a trav�s de D1 y D2.
�   '    �  -����Arial����                       Arial            
 #�@ ����        ��������#�             0     ��������#� ����      @5     ��������#�  ʚ;�������?.1     ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true
     ��������#� ����  false     ��������               
                  #� ����        ��������#� ����       ��������#�  ����       ��������#�@ ����       ��������#�@ ����       ��������               
                  #� ����        ��������#� ����       ��������#�@ ����       ��������#�  ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������               
                 #� ����dec     ��������#� ����     @�@1k     ��������#� ����    ��.A1meg     ��������#� ����       20     ��������#� ���� true     ��������#� ���� true     ��������#� ���� true	     ��������#� ����  false
     ��������               
                 #�  ����        ��������#�  ����       ��������#�  ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������               
                  	 #� ����        ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������               
                 #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
                    #�             0      ��������#�  ��{�G�z�?20m     ��������#�  � -C��6
?0.05m     ��������#�  � -C��6
?0.05m     ��������#� ���� True     ��������#� ����  F     ��������#� ���� true     ��������#� ����  false     ��������               
                 #� ����     @�@1K      ��������#�  ����       ��������#�  ����       ��������#�  ����       ��������               
         ��              #�  ����        ��������              
                  #�  ����        ��������              
                                  
                 #�@ ����        ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true	     ��������#� ����  false
     ��������#� ���� true     ��������#� ����  false     ��������               
                 #� ����       5      ��������#� ����       5     ��������#� ����       5     ��������#� ����       5     ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#�@ ����       ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#� ���� true     ��������#� ���� true     ��������#� ����  false     ��������#� ���� true     ��������#� ����  false      ��������#� ���� true!     ��������#� ����  false"     ��������               
                        #� ����       5      ��������#� ����       5     ��������#� ����       5     ��������#� ����       5     ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#�@ ����       ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#� ���� true     ��������#� ���� true     ��������#� ����  false     ��������#� ���� true     ��������#� ����  false      ��������#� ���� true!     ��������#� ����  false"     ��������               
                 #� ����       5      ��������#� ����       5     ��������#� ����       5     ��������#� ����       5     ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#�@ ����       ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#� ���� true     ��������#� ���� true     ��������#� ����  false     ��������#� ���� true     ��������#� ����  false      ��������#� ���� true!     ��������#� ����  false"     ��������               
                 #� ����       5      ��������#� ����       5     ��������#� ����       5     ��������#� ����       5     ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#�@ ����       ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#� ���� true     ��������#� ���� true     ��������#� ����  false     ��������#� ���� true     ��������#� ����  false      ��������#� ���� true!     ��������#� ����  false"     ��������               
                 #�@ ����        ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����decade     ��������#� ���� true     ��������#� ���� true     ��������#� ���� true     ��������#� ����  false     ��������               
                 #� ����        ��������#� ����       ��������#�@ ����       ��������#�  ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������               
                        #� ����dec     ��������#� ����     @�@1k     ��������#� ����    ��.A1meg     ��������#� ����       20     ��������#� ����        0     ��������#� ����        0     ��������#� ���� true	     ��������#� ���� true
     ��������#� ����      I@50     ��������#� ���� true     ��������#� ����  false     ��������               
                         / #� ���� x'     ��������#�     �-���q=1E-12     ��������#� @B -C��6?1E-4     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x	     ��������#� ���� x!     ��������#� ����    �  500
     ��������#� ���� x     ��������#� ����    �  500     ��������#� ���� x$     ��������#� ���� x$     ��������#� ���� x%     ��������#� ���� x"     ��������#�  ���� x*     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x&     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x+     ��������#� ���� x,     ��������#� ���� x-     ��������#� ���� xg     ��������#� ���� xf     ��������#� ���� xd     ��������#� ���� xe     ��������#� ���� xh     ��������#� ���� xj     ��������#� ���� xi     ��������#� ���� xk     ��������#� ����    e��A1Gl     ��������#�             0�     ��������#� ����      @5�     ��������#� ����      @2.5�     ��������#� ����      �?.5�     ��������#� ����      @4.5�     ��������#� 
   ��&�.>1n�     ��������#� 
   ��&�.>1n�     ��������#� 
   ��&�.>1n�     ��������#� 
   ��&�.>1n�     ��������           ��  CPrimitiveModel    d1n4007   #�    1�a��%>2.55e-9      ��������#� ���� 27     ��������#�  �/�$��?0.042     ��������#� ����      �?1.75     ��������#�  �  ��v��(�>5.76e-6     ��������#�     �]}IW�=1.85e-11     ��������#� ����      �?0.75     ��������#� ����Zd;�O�?0.333     ��������#� ���� 1.11	     ��������#� ���� 3.0
     ��������#�      0     ��������#� ���� 1     ��������#� ���� 0.5     ��������#� ����     @�@1000     ��������#� � Ǯ���?9.86e-5     ��������     Diode Generic��   CPrimitiveModelType Junction Diode model����DD   >����� 1.0E-14Saturation current    ProcessisAmp0       e     >����� 27!Parameter measurement temperature    ProcesstnomDeg C0     s     >����� 0Ohmic resistance    ProcessrsOhm0      f     >����� 1Emission Coefficient    Processn 0      g     >����� 0Transit Time    Processttsec0     h     >����� 0Junction capacitance    ProcesscjoF0     i     >����� 0     Processcj0F0     i     >����� 1Junction potential    ProcessvjV0      j     >����� 0.5Grading coefficient    Processm 0      k     >����� 1.11Activation energy    ProcessegeV0     	 l     >����� 3.0#Saturation current temperature exp.    Processxti 0     
 m     >����� 0flicker noise coefficient    Processkf 0      t     >����� 1flicker noise exponent    Processaf 0      u     >����� 0.5#Forward bias junction fit parameter    Processfc 0      n     >����� infReverse breakdown voltage    ProcessbvV0      o     >����� 1.0e-3$Current at reverse breakdown voltage    ProcessibvA0      p     >�����  Ohmic conductance    ProcesscondMho     r        D��     9I�                Ariald         �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ ��  COpAnal                         
                        ����            
H13               ��  TSignal                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                      v(iv_vl)       ����                  ʃ                     	i(va_ix1)       ����                  ʃ                     i(itiristor)       ����                  ʃ                     i(va_il)       ����                  ʃ                      	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ ��  CDCsweep       
 ����������               
                       ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                       v(iv_vl)       ����                  ʃ                      	i(va_ix1)       ����                  ʃ                      i(itiristor)       ����                  ʃ                      i(va_il)       ����                  ʃ                       	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ ��  CACsweep        ��������               
                       ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                      v(iv_vl)       ����                  ʃ                     	i(va_ix1)       ����                  ʃ                     i(itiristor)       ����                  ʃ                     i(va_il)       ����                  ʃ                      	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ �� 
 CTranSweep       ��������               
                       ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                       v(iv_vl)       ����                  ʃ                      	i(va_ix1)       ����                  ʃ                      i(itiristor)       ����                  ʃ                      i(va_il)       ����                  ʃ                       	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ ��  CACdisto        �����               
                           ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                       v(iv_vl)       ����                  ʃ                      	i(va_ix1)       ����                  ʃ                      i(itiristor)       ����                  ʃ                      i(va_il)       ����                  ʃ                       	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ �        #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
         �                 ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                       v(iv_vl)       ����                  ʃ                      	i(va_ix1)       ����                  ʃ                      i(itiristor)       ����                  ʃ                      i(va_il)       ����                  ʃ                       	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ �        #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
         �                 ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                       v(iv_vl)       ����                  ʃ                      	i(va_ix1)       ����                  ʃ                      i(itiristor)       ����                  ʃ                      i(va_il)       ����                  ʃ                       	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ �        #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
         �                 ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                       v(iv_vl)       ����                  ʃ                      	i(va_ix1)       ����                  ʃ                      i(itiristor)       ����                  ʃ                      i(va_il)       ����                  ʃ                       	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ �        #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
         �                 ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                       v(iv_vl)       ����                  ʃ                      	i(va_ix1)       ����                  ʃ                      i(itiristor)       ����                  ʃ                      i(va_il)       ����                  ʃ                       	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ �        #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
         0             	    ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                      v(iv_vl)       ����                  ʃ                     	i(va_ix1)       ����                  ʃ                     i(itiristor)       ����                  ʃ                     i(va_il)       ����                  ʃ                      	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ ��  CACnoise        ��������               
                    
    ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                      v(iv_vl)       ����                  ʃ                     	i(va_ix1)       ����                  ʃ                     i(itiristor)       ����                  ʃ                     i(va_il)       ����                  ʃ                      	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ ��         #�  ����        ��������#�  ����       ��������#�  ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������              
                        ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                      v(iv_vl)       ����                  ʃ                     	i(va_ix1)       ����                  ʃ                     i(itiristor)       ����                  ʃ                     i(va_il)       ����                  ʃ                      	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ ��  CFourier        ����               
         ��                   ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                      v(iv_vl)       ����                  ʃ                     	i(va_ix1)       ����                  ʃ                     i(itiristor)       ����                  ʃ                     i(va_il)       ����                  ʃ                      	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ ��  CACpz        	 ���������               
                       ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                      v(iv_vl)       ����                  ʃ                     	i(va_ix1)       ����                  ʃ                     i(itiristor)       ����                  ʃ                     i(va_il)       ����                  ʃ                      	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ ��  CDCtf         �����               
                       ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                      v(iv_vl)       ����                  ʃ                     	i(va_ix1)       ����                  ʃ                     i(itiristor)       ����                  ʃ                     i(va_il)       ����                  ʃ                      	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ ��  CDCsens         �����������               
                       ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                       v(iv_vl)       ����                  ʃ                      	i(va_ix1)       ����                  ʃ                      i(itiristor)       ����                  ʃ                      i(va_il)       ����                  ʃ                       	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ                 ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                      v(iv_vl)       ����                  ʃ                     	i(va_ix1)       ����                  ʃ                     i(itiristor)       ����                  ʃ                     i(va_il)       ����                  ʃ                      	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ ��  CShow         �              
                       ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                      v(iv_vl)       ����                  ʃ                     	i(va_ix1)       ����                  ʃ                     i(itiristor)       ����                  ʃ                     i(va_il)       ����                  ʃ                      	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ ��  CShowmod         �              
                       ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                      v(iv_vl)       ����                  ʃ                     	i(va_ix1)       ����                  ʃ                     i(itiristor)       ����                  ʃ                     i(va_il)       ����                  ʃ                      	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ �� 
 CLinearize        #�  ����        ��������               
                       ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                      v(iv_vl)       ����                  ʃ                     	i(va_ix1)       ����                  ʃ                     i(itiristor)       ����                  ʃ                     i(va_il)       ����                  ʃ                      	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ ��  CParamTranSweep        �������������               
                       ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                      v(iv_vl)       ����                  ʃ                     	i(va_ix1)       ����                  ʃ                     i(itiristor)       ����                  ʃ                     i(va_il)       ����                  ʃ                      	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ �              ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                       v(iv_vl)       ����                  ʃ                      	i(va_ix1)       ����                  ʃ                      i(itiristor)       ����                  ʃ                      i(va_il)       ����                  ʃ                       	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ ��  CParamACSweep        RSTUVWXYZ[\]^               
                       ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                      v(iv_vl)       ����                  ʃ                     	i(va_ix1)       ����                  ʃ                     i(itiristor)       ����                  ʃ                     i(va_il)       ����                  ʃ                      	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ ��  CMonteCarlo_op        ����������������������������               
                              ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                      v(iv_vl)       ����                  ʃ                     	i(va_ix1)       ����                  ʃ                     i(itiristor)       ����                  ʃ                     i(va_il)       ����                  ʃ                      	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ ��  CMonteCarlo_dc        �� 	
               
                       ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                       v(iv_vl)       ����                  ʃ                      	i(va_ix1)       ����                  ʃ                      i(itiristor)       ����                  ʃ                      i(va_il)       ����                  ʃ                       	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ ��  CMonteCarlo_ac         !"#$%&'()*+,-./012345               
                       ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                      v(iv_vl)       ����                  ʃ                     	i(va_ix1)       ����                  ʃ                     i(itiristor)       ����                  ʃ                     i(va_il)       ����                  ʃ                      	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ ��  CMonteCarlo_tran        6789:;<=>?@ABCDEFGHIJKLMNOPQ               
                       ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                       v(iv_vl)       ����                  ʃ                      	i(va_ix1)       ����                  ʃ                      i(itiristor)       ����                  ʃ                      i(va_il)       ����                  ʃ                       	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ ��  CACsens        _`abcdefghi               
                              ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                       v(iv_vl)       ����                  ʃ                      	i(va_ix1)       ����                  ʃ                      i(itiristor)       ����                  ʃ                      i(va_il)       ����                  ʃ                       	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ ��  CNetworkAnalysis        jklmnopqrst               
                       ����            P               ʃ                        v(ctrl)       ����                  ʃ                       v(13)       ����                  ʃ                       v(3)       ����                  ʃ                       v(4)       ����                  ʃ                       v(5)       ����                  ʃ                       v(9)       ����                  ʃ                       v(6)       ����                  ʃ                       v(11)       ����                  ʃ                       v(10)       ����                  ʃ	                       i(v1)       ����                  ʃ
                       v(iv_vl)       ����                  ʃ                      	i(va_ix1)       ����                  ʃ                      i(itiristor)       ����                  ʃ                      i(va_il)       ����                  ʃ                       	v(iv_vx1)       ����                      �O�{��3 ��3 t�3 v�{�6ϑ     �O�{��3 ��3 t�3 v�{�6ϑ                 ����            P                 >           ��   CDigSimResTemplate                ���       ����  ����:�0�yU>20.00n���   ����                       Arial����                       Arial����                       Arial  �   �  �                                ����  ���� ������       ����  ���� ������                 �               ����  �����       200������         0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial      �       �         �     �   �  �  Circuit1                  ����  ��    ��������                                                                                                                                                                                                                           g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     ��   CPackageAliasSuperPCBStandardDIODE3      ЅEagle	DIODE.LBRDO41-7   AC  ЅOrcad 	DAX2/DO41      Ѕ	Ultiboard	L7DIO.l55DIO_DO41              A      g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     ЅSuperPCBStandardDIODE3      ЅEagle	DIODE.LBRDO41-7   AC  ЅOrcad 	DAX2/DO41      Ѕ	Ultiboard	L7DIO.l55DIO_DO41              A                                                �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                     CM�� ����P�3     ��3 ���{                      .:\�`�              2         �  �              � � �           ��3     ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                      �                  ��         �  @                  ���                                                  �  @  �     <   �  <     ��                                                        �     |   �  |     ��                                                        �     �   �  �     ��                                                        �     �   �  �     ��                                                        � �      �  4     ��                                                      �      �  4   �      �  4   [title]                                       � �   D   �  t     ��                                                      �   D   �  t   �   D   �  t   [description]                                       � `   �   h  �     ��                                                      `   �   h  �   `   �   h  �   [id]                                       � �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       �      �   8    ��        	                                                   �   8       �   8  Date :       �  ,  H  �                  � �     �  4   	 ��        
                                              �     �  4  �     �  4  [date]                                       �       t   8    
 ��                                                            t   8         t   8   Title :       �  ,     �                  �    L   �   x     ��                                                         L   �   x      L   �   x   Description :       �  �  �   �                  �    �   �   �     ��                                                         �   �   �      �   �   �   ID :       �  �  �  V                  �    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �  l  8                      ��������������          �     	title box    Analog Misc      �?    9 
 8�     #�  ����        ��������#�  ����       ��������#�  ����       ��������#�  ����       ��������#�  ����       ��������        9                                      ����<��� ����     >�            title                >�            description               >�            id               >�            designer               >�            date                           ����            `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                                                                                            2         �  �              � � �                   ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                          �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   
cgs 76         47 80moh5.6 L2 �S��
mvrd nmodel `�w    37     ʃ                      TIME� # ) time                      ʃ                        i(v1)� < � i(v1)    TIME                 ʃ                        v(3)      v(3)    TIME                 ʃ                      	i(va_ix1)�   � 	i(va_ix1)    TIME                 ʃ    (v(7)-v(3))                   v(IV_VL)� �   v(IV_VL)    TIME                 ʃ                      i(va_il)  � � i(va_il)    TIME                 ʃ    v(5)                   	v(IV_Vx1)� �   	v(IV_Vx1)    TIME                 ʃ    v(iv_vx1)*i(va_ix1)                    Pin� # )  ����TIME                 ʃ                        v(ctrl)      v(ctrl)    TIME                 ʃ                        v(5)      v(5)    TIME                 ʃ                        v(ctrl2)      v(ctrl2)    TIME                           2         �  �           Time  � � �             �?    ����                       Arial����                       Arial                              ����  �����z�`?2.035181e-003��G�6      ����  �����z�`?2.035181e-003��G�6      ����  ����1��{��%�-1.075922e+001������      ����  ����1��{��%�-1.075922e+001������                                                                         �                      �                                                                                                                                                                                                                                                                                                                                                                                          �  �                                                                                                                                                                                                                                                                                                                                                                                                  �  �                                              �                      �                              1m  0                            100   100                                                             1m  0                            100   100                                1m  0                            100   100                                1m  0                            100   100                                                 
                 1m  0                            100   100                            ��   CPartPackage     ��   CPackageg   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     ����   ��/� �g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     ����      ��   CMiniPartPin    ����V+V+     PWR+V+g      	�   ����V-V-     PWR-V-h     voltage_sourcevoltage_source                          	�    ����C+C+     PASC+�      	�   ����C-C-     PASC-�     capacitor_genericcapacitor_generic                          	�    ����11     PAS1�      	�   ����22     PAS2�     BatteryBattery                          	�    ����R+R+     PASR+      	�   ����R-R-     PASR-     RR                          	�    ����GndGnd     GNDGnd}      GndGnd                  	�    ����M+M+     PASM+i      	�   ����M-M-     PASM-j     	voltmeter	voltmeter                          	�    ����M+M+     PASM+2      	�   ����M-M-     PASM-3     Ammeter2Ammeter2                          	�    ����MM       ��������MarkerMarker                  	�    ����GndGnd     GNDGnd}      GndGnd                  	�    ����GndGnd     GNDGnd}      GndGnd                  	�    ����11     PAS1S      	�   ����22     PAS2T     	�   ����33     PAS3U     	�   ����44     PAS4V     vcswitchvcswitch                                          	�    ����GndGnd     GNDGnd}      GndGnd                  	�    ����MM       ��������MarkerMarker                  	�    ����L+L+     PASL+K      	�   ����L-L-     PASL-L     InductorInductor                          	�    ����M+M+     PASM+0      	�   ����M-M-     PASM-1     AmmeterAmmeter                          	�    ����M+M+     PASM+k      	�   ����M-M-     PASM-l     
Voltmeter2
Voltmeter2                        	�    ����D+D+     PASA       	�   ����D-D-     PASK       �   ��   CPackagePin 1 D+PAS  AA(� 2 D-PAS  AKDiodeDiode	Fairchild      1n4007 D1n4007D2            diode-21n40071n4007                        	�    ����D+D+     PASA       	�   ����D-D-     PASK       C  (� 1 D+PAS  AA(� 2 D-PAS  AKDiodeDiode	Fairchild      1n4007 D1n4007D1            diode-21n40071n4007                          	�    ����GndGnd     GNDGnd}      GndGnd                  	�    ����11     PAS1S      	�   ����22     PAS2T     	�   ����33     PAS3U     	�   ����44     PAS4V     vcswitchvcswitch                                          	�    ����V+V+     PWR+V+g      	�   ����V-V-     PWR-V-h     voltage_sourcevoltage_source                                                                                                                                                                                         
m1     8 8 mm l=100u w                        used                            ��    �Z�P��,�                        ��                                                                                                            (f    x=f � �'f                           �(f                            ,�e    �f � ��e                           ��e                                     �  � ���� �                         .I                                                                                                                                                                                                                                                                                                                                                       �$�    h&��&��&� '�                        H)�                            MJ         W X Y [   Z                          DIN                            sist      resistor DIN                                                       ��    ��������P��                        ��                            �V�    (W�`W��W��W�                        �Y�                            Їl    `�l(�l`-j �W                         �W                            t�@
    L �k��
>ENDDATA
                        
JV1                            p�<        ��<x�                           �                                         �rP��                                                                                                                                                      �rP��                                 2 2 2 2 d                                                                               