    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz        ��  CPart           �   �          �   �              Battery��  CIntPin    ��  CWire     �      �	       �      �      �      �              ua555�         4 �   �    �       �       _      �      _      �              capacitor_generic �   �     �         �           �   �           �   �               Gnd ��  CExtPin    ��  CVertex   �  �
   ��  CSegment   �   �                    �,    �&   �  �
   �    �   �   
                   �+    �;    	  �
   �3   �    	  �        	                                        `       Gnd}   @  �
          gnd1     ��   CPin                    ��                                                               Gnd��  TLine                   ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        #�         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        #�    ,   4   ,     ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        #�    8   (   8     ��    p�Z         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         " $ % '   &      Ground    
Ground DINMiscellaneous      �?       ��   CGroundBehavior       Gnd ��   CBehPin     Gnd        ����Gnd����                        ��gndgnd                 + Analog Meters   Generic   gnd1gnd1          ����  gnd ��   CPartPin    ����GndGnd      GNDAGnd    ����SourcesGroundGeneric              0 �        0  �        0  *�    2      ����2����                        ��+ *�    C-      ����C-����                        ��*�    ground����   ����GROUND����                        ��  0     0 �           �  C-�  �   �    �  @   �7   5 �A   �  �   6 �/   �    �      �2   �?   �  `   : �.   ; �	   �  `   <                9     8 �(   9 �0          >    	            7     �*   7 �      �   @    	                              �   C+�   �  �         C     !�                   ��                                                           �   C-!�                   ��                                                          @   C+#�     @       �      ��    
*                                                 #�     �   �����     ��     gro                                                #�     �   �����     ��     
q                                                #�     �       �     ��    jt_n                                                ��  
 TTextField 0   t   �   �     ��                                                       0   t   �   �   0   t   �   �   [capacitance]         �  �  r	      `   �   �   H� 0   @   �   d     ��                                                       0   @   �   d   0   @   �   d   	[refname]         @  X  �          �   $    D E F G I     J       B C  �  	Capacitor     Miscellaneous      �?       ��  CCapacitorBehavior     ��  CValue '  Vo�c�/4>4.7n      ��������M� ���� x     ��������M� ����       ��������M� ����       �������� C+C- *�     C+        ����C+����                        ��1  	capacitor   i            R 1 Passive   Generic   CC          ����  C ,�    ����C+C+      PASAC+��X����,�   ����C-C-      PASAC-�<
����Passive Generic              3 �      �       �   �  �       �   �  �               resistor_generic�    �    �    X    �   /   �      �   /   �      �               MarkerY �    �<    
  `   �1   �    	  `   ]    	    \     �0   �>    
  `   �6   �
   @  `   a         `     _     \                `      M     �	  @         Vout     !�                   ��                                                           `   M#� 0   `       `     ��    ���                                                 ��  TPolygon �����  �����     ��                                                         ��  TPointP   `    pQg�@   P       g�0   `        g�@   p            H� `   P      t     ��                                                       `   P      t   `   P      t   	[refname]       �
  0  �  �        �   ,    f   c l d  �  Marker     Miscellaneous      �?    +   ��   CMarkerBehavior     M�             0.0      �������� M ��  	 TModelPin ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     X n   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               q Analog MiscV   Generic   VoutVout          ����               Vout  v(Vout)  N ,�    ����MM       A    ����RootmarkerGeneric              Vout �   X    Vout W  *�     R+        ����R+����                        ��*�    out����   ����out����                        ��q  Vout   V Vout U �    b    �  �   R+  �   =       �   R-   �  �         RA     !�                    ��                                                       �   @   R+!�                   ��                                                          @   R-#�    @   $   0     ��    �                                                 #� 0   P   $   0     ��                                                       #� 0   P   <   0     ��    ��K                                                #� H   P   <   0     ��                                                       #� H   P   T   0     ��                                                        #� `   P   h   @     ��    (�K                                                #� �   @   h   @     ��                                                       #� `   P   T   0    	 ��        	                                                #�    @       @    
 ��        
                                                H�     `   �   �     ��                                                           `   �   �       `   �   �   [resistance]       �  �  (  V      `   �   �   H�         t   $     ��                                                               t   $           t   $   	[refname]       �  �  P  @          t   $    x y z { | } ~  � � � � �    resistor    resistor DINMiscellaneous      �?       ��  CResistorBehavior     M� ����     @�@2k      ��������M� ���� 27     ��������M� ����       ��������M� ����       �������� R+R- t *�    R-      ����R-����                        �� resistor   i            t � Passive   Generic   RARA          ����    R ,�    ����R+R+      PASAR+G3 ����,�   ����R-R-      PASAR-DATA����Passive Generic              3 
 �       3  R � *�    thr����   ����thr����                        ��*�    trg����   ����trg����                        �� 3   3 �   �    �  *�    ctrl����   ����ctrl����                        �� 5   5 �  �   �    �  *�    dis����   ����dis����                        �� 2   2 s / �    �!      �   �)   �   �  �   �4   � �@   �  �   � �-   � �=    	  �   �5   � �    	  �   �    	        �                 �         �        	               VCC:  �   ?       �  	THRESHOLD;  �   �      `       	          �  Control<  �   A       @  TRIGGER=  �   �         RESET>  �   �    	          	         �  	DISCHARGE?  �   ^      �  OUTPUT@  �          @  GROUNDA      �          U1     !�                    ��                                                           `   VCC!�                   ��                                                          �   	THRESHOLD!�                   ��                                                          �   Control!�                   ��                                                          �   TRIGGER!�                   ��                                                         `   RESET!�                   ��                                                         �   	DISCHARGE!�                   ��                                                         �   OUTPUT!�                   ��                                                         �   GROUND#�     `       `    	 ��                                                        #�     �       �    
 ��        	                                                #�     �       �     ��        
                                                #�     �       �     ��                                                        #� �   `      `     ��                                                        #� �   �      �     ��     ��                                                #� �   �      �     ��                                                        #� �   �      �     ��     �                                                 �� 
 TRectangle     @   �   �                  ����                                             @   �   �   H� (   P   p   p     ��                                                      (   P   p   p   (   P   p   p   vcc       x  p  �  �  (   P   p   p   H� (   p   p   �     ��                                                      (   p   p   �   (   p   p   �   thr       x  �  �  R  (   p   p   �   H� (   �   p   �     ��                                                      (   �   p   �   (   �   p   �   cont       x  0    �  (   �   p   �   H� (   �   p   �     ��                                                      (   �   p   �   (   �   p   �   trIg       x  �  �    (   �   p   �   H� �   P   �   p     ��                                                      �   P   �   p   �   P   �   p   reset       �  p  H  �  �   P   �   p   H� �   p   �   �     ��                                                      �   p   �   �   �   p   �   �   dischg       �  �  �  R  �   p   �   �   H� �   �   �   �     ��                                                      �   �   �   �   �   �   �   �   out       �  0    �  �   �   �   �   H� �   �   �   �     ��                                                      �   �   �   �   �   �   �   �   gnd       �  �  (    �   �   �   �   H�     �����        ��                                                           �����          �����      	[devname]        ����������������    �����      H�        �   <     ��                                                              �   <          �   <   	[refname]       `  �  �  h         �   <    � � � � � � � � �   � � � � � � � � � � � � � � � � � �      lm555     Miscellaneous      �?   #    U ,�    ����VCCvcc      PASAVCC    ����,�   ����	THRESHOLDthr      PASA	THRESHOLD    ����,�   ����Controlctrl      PASAControl    ����,�   ����TRIGGERtrg      PASATRIGGER4   ����,�   ����RESETrst      PASARESET   �����,�   ����	DISCHARGEdis      PASA	DISCHARGE0'3����,�   ����OUTPUTout      PASAOUTPUT    ����,�   ����GROUNDground      PASAGROUND��Z����Timer	555 timerNational Semiconductor              4 	  *�     1       ����1����                        ��*�     vcc����    ����vcc����                        ��*�    rst����   ����rst����                        �� 4    4 . �    �    `       1�  �      `   �  2�   @  �          X1     !�                    ��                                                               1!�                   ��                                                          �   2#�             $     ��    ��)                                                #�     \       �     ��                                                        #�    8   0   8    	 ��    ��)                                                #�     H   @   H     ��    p�Z                                                #�     $   @   $     ��                                                       #�    \   0   \     ��    D�Z                                                #�               ���                                                      #�               ���   �Z	                                                H� `          $    
 ��        
                                               `          $   `          $   	[devname]        ����������������`          $   H� `   $      H     ��                                                       `   $      H   `   $      H   	[refname]       `    �  �  `   $      H    � � � � � � � �     � �     �   �      Battery     Miscellaneous      �?    9 
 ��  CParamSubBehavior     M� ����      (@12      �������� 12 � 0 BatteryBattery  9 i             � 0 Sources   Generic   X1X1          ������   CParamSubModelType��    BATTERY2.SUBCKT Xbattery 1 2
V1 1 2 DC {voltage}
.ENDS
   ��  	 CParmDefn    1battery voltage   ParamSubvoltageV                X ,�    ����11      PASA1�1b����,�   ����22      PASA2�Y����SourcesBatteryGeneric                  V                  Z     X   � � 8  8                                                                               > � @   � < 8 _ ] :  � � a 6 B  B 5               = b �           �                  ^   � A � 9 �                            ?                      \ � ` ; � 7    ��  CLetter    T = 1.76 * RA * C  _  �  �      ����Arial����                       Arial     �   =Ajustant Ra i C, podem ajustar la frencuencia de l'oscilador.w  /  H  �      ����Arial����                       Arial     �   �6C           R              T                F
4.7n      250         2 us          480 kHz
4.7n      500        4.1 us        240 kHz
4.7n       1k         8.2 us        120 kHz
4.7n       2k        16.4 us        60 kHz
4.7n       10k        82 us         12 kHz
4.7n       20k       164 us         6 kHzw  �    �      ����Arial����                       Arial     �   �Substituint RA per una resistencia de 250 ohms en serie
amb un potenci�metre de 20 kohms ens ha de permetre
modificar la frencuencia de 555 de 5 kHz a 500 kHz aprox.�  �  �  �      ����Arial����                       Arial            
 M�@ ����        ��������M�             0     ��������M� ����      @5     ��������M�  ʚ;�������?.1     ��������M�@ ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ���� true
     ��������M� ����  false     ��������               
                  M� ����        ��������M� ����       ��������M�  ����       ��������M�@ ����       ��������M�@ ����       ��������               
                  M� ����        ��������M� ����       ��������M�@ ����       ��������M�  ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������               
                 M� ����dec     ��������M� ����     @�@1k     ��������M� ����    ��.A1meg     ��������M� ����       20     ��������M� ���� true     ��������M� ���� true     ��������M� ���� true	     ��������M� ����  false
     ��������               
                 M�  ����        ��������M�  ����       ��������M�  ����       ��������M� ����dec     ��������M� ����       ��������M� ����       ��������M� ����  	     ��������M� ����  
     ��������               
                  	 M� ����        ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������               
                 M� ����        ��������M� ����       ��������M� ����       ��������M� ����dec     ��������M� ����       ��������               
                    M�             0      ��������M� @B ,C��6?100u     ��������M� �  H�����z>0.1u     ��������M� �  H�����z>0.1u     ��������M� ���� True     ��������M� ����  F     ��������M� ���� true     ��������M� ����  false     ��������               
                 M� ����     @�@1K      ��������M�  ����       ��������M�  ����       ��������M�  ����       ��������               
         ��              M�  ����        ��������              
                  M�  ����        ��������              
                                  
                 M�@ ����        ��������M�@ ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ���� true	     ��������M� ����  false
     ��������M� ���� true     ��������M� ����  false     ��������               
                 M� ����       5      ��������M� ����       5     ��������M� ����       5     ��������M� ����       5     ��������M� ����       ��������M� ����  	     ��������M� ����  
     ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ���� true     ��������M�@ ����       ��������M�@ ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����dec     ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ���� true     ��������M� ���� true     ��������M� ���� true     ��������M� ����  false     ��������M� ���� true     ��������M� ����  false      ��������M� ���� true!     ��������M� ����  false"     ��������               
                        M� ����       5      ��������M� ����       5     ��������M� ����       5     ��������M� ����       5     ��������M� ����       ��������M� ����  	     ��������M� ����  
     ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ���� true     ��������M�@ ����       ��������M�@ ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����dec     ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ���� true     ��������M� ���� true     ��������M� ���� true     ��������M� ����  false     ��������M� ���� true     ��������M� ����  false      ��������M� ���� true!     ��������M� ����  false"     ��������               
                 M� ����       5      ��������M� ����       5     ��������M� ����       5     ��������M� ����       5     ��������M� ����       ��������M� ����  	     ��������M� ����  
     ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ���� true     ��������M�@ ����       ��������M�@ ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����dec     ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ���� true     ��������M� ���� true     ��������M� ���� true     ��������M� ����  false     ��������M� ���� true     ��������M� ����  false      ��������M� ���� true!     ��������M� ����  false"     ��������               
                 M� ����       5      ��������M� ����       5     ��������M� ����       5     ��������M� ����       5     ��������M� ����       ��������M� ����  	     ��������M� ����  
     ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ���� true     ��������M�@ ����       ��������M�@ ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����dec     ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ���� true     ��������M� ���� true     ��������M� ���� true     ��������M� ����  false     ��������M� ���� true     ��������M� ����  false      ��������M� ���� true!     ��������M� ����  false"     ��������               
                 M�@ ����        ��������M�@ ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����decade     ��������M� ���� true     ��������M� ���� true     ��������M� ���� true     ��������M� ����  false     ��������               
                 M� ����        ��������M� ����       ��������M�@ ����       ��������M�  ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������M� ����       ��������               
                        M� ����dec     ��������M� ����     @�@1k     ��������M� ����    ��.A1meg     ��������M� ����       20     ��������M� ����        0     ��������M� ����        0     ��������M� ���� true	     ��������M� ���� true
     ��������M� ����      I@50     ��������M� ���� true     ��������M� ����  false     ��������               
                         / M� ���� x'     ��������M�     �-���q=1E-12     ��������M� @B -C��6?1E-4     ��������M� ���� x     ��������M� ���� x     ��������M� ���� x     ��������M� ���� x     ��������M� ���� x     ��������M� ���� x     ��������M� ���� x	     ��������M� ���� x!     ��������M� ����    �  500
     ��������M� ���� x     ��������M� ����    �  500     ��������M� ���� x$     ��������M� ���� x$     ��������M� ���� x%     ��������M� ���� x"     ��������M�  ���� x*     ��������M� ���� x     ��������M� ���� x     ��������M� ���� x     ��������M� ���� x&     ��������M� ���� x     ��������M� ���� x     ��������M� ���� x     ��������M� ���� x+     ��������M� ���� x,     ��������M� ���� x-     ��������M� ���� xg     ��������M� ���� xf     ��������M� ���� xd     ��������M� ���� xe     ��������M� ���� xh     ��������M� ���� xj     ��������M� ���� xi     ��������M� ���� xk     ��������M� ����    e��A1Gl     ��������M�             0�     ��������M� ����      @5�     ��������M� ����      @2.5�     ��������M� ����      �?.5�     ��������M� ����      @4.5�     ��������M� 
   ��&�.>1n�     ��������M� 
   ��&�.>1n�     ��������M� 
   ��&�.>1n�     ��������M� 
   ��&�.>1n�     ��������                 � ��  CMacroBehavior      vccthrctrltrgrstdisoutground � � � � � � u 2 ua555ua555 # u             � � � � � � u 2 Timer�   Generic   U1U1          ��************************
* B2 Spice Subcircuit
************************
* Pin #		Pin Name
* vcc		vcc
* thr		thr
* ctrl		ctrl
* trg		trg
* rst		rst
* dis		dis
* out		out
* GROUND		GROUND
.Subckt ua555 vcc thr ctrl trg rst dis out GROUND 


***** main circuit
R1 vcc  9  4.7K 
R2 vcc  3  830 
R3 vcc  8  4.7k 
R4 vcc  10  1K 
R5 vcc  ctrl  5K 
R7 17  0  10K 
Q6 2  thr  5 bjt_npn_generic 
Q2 25  2  3 bjt_pnp_generic 
Q3_ 0  6  3 bjt_pnp_generic 
Q1 2  2  9 bjt_pnp_generic 
Q7 2  5  17 bjt_npn_generic 
Q8 6  4  17 bjt_npn_generic 
Q9 6  ctrl  4 bjt_npn_generic 
Q4 6  6  8 bjt_pnp_generic 
Q5 12  20  10 bjt_pnp_generic 
Q17_ 15  rst  31 bjt_pnp_generic 
Q16 dis  15  0 bjt_npn_generic 
R14_ 15  16  100 
Q14_ 0  trg  11 bjt_pnp_generic 
Q12_ 22  11  12 bjt_pnp_generic 
Q13_ 14  13  12 bjt_pnp_generic 
Q15_ 14  18  13 bjt_pnp_generic 
R8_ 22  0  100K 
R0 ctrl  18  5K 
R10 18  0  5K 
Q21_ 25  22  0 bjt_npn_generic 
Q20_ 24  25  0 bjt_npn_generic 
Q22_ 27  24  0 bjt_npn_generic 
Q24_ 29  27  16 bjt_npn_generic 
Q25_ out  26  0 bjt_npn_generic 
Q23_ vcc  29  28 bjt_npn_generic 
Q26 vcc  28  out bjt_npn_generic 
Q19 20  20  vcc bjt_pnp_generic 
R11_ 20  31  5K 
D1 31  24 diode 
R12_ 25  27  4.7K 
R15_ 16  26  220 
R16_ 16  0  4.7K 
D2 out  29 diode 
R6_ vcc  29  6.8K 
R17_ 28  out  3.9K 
R9_ 14  0  100K 
Q18 27  20  vcc bjt_pnp_generic 

.model bjt_npn_generic npn  is = 5f   bf = 100    nf = 1   vaf = 160   ikf = 30m   ise = 4p  
+ ne = 2   br = 4   nr = 1   var = 16   ikr = 45m  
+ rb = 4   re = 1.0   rc = .4   cje = 12.4p   vje = 1.1  
+ mje = .5   tf = 250p   cjc = 4p   vjc = .3   mjc = .3  
+ tr = 1n  

.model bjt_pnp_generic pnp  is = 1.0e-14   bf = 20    vaf = 50   ne = 2   br = .02   rb = 25  
+ rc = 4   cje = 12.4p   vje = 1.1   mje = .5   tf = 250p  
+ vjc = .3   mjc = .3   tr = 100n  

.model diode D  is = 1.0E-14   rs = 40   cjo = 1p  

.ends                 Ariald     ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j                   ����            > A               ��  TSignal                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  ��  CDCsweep       
 � � � � � � � � � �                
                       ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  ��  CACsweep        	
               
                       ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  �� 
 CTranSweep       %&'()*+,               
                       ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  ��  CACdisto         !"#$               
                           ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  �        M� ����        ��������M� ����       ��������M� ����       ��������M� ����dec     ��������M� ����       ��������               
         �                 ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  �        M� ����        ��������M� ����       ��������M� ����       ��������M� ����dec     ��������M� ����       ��������               
         �                 ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  �        M� ����        ��������M� ����       ��������M� ����       ��������M� ����dec     ��������M� ����       ��������               
                           ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  �        M� ����        ��������M� ����       ��������M� ����       ��������M� ����dec     ��������M� ����       ��������               
         �                 ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  �        M� ����        ��������M� ����       ��������M� ����       ��������M� ����dec     ��������M� ����       ��������               
                      	    ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  ��  CACnoise                       
                    
    ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  ]�         M�  ����        ��������M�  ����       ��������M�  ����       ��������M� ����dec     ��������M� ����       ��������M� ����       ��������M� ����  	     ��������M� ����  
     ��������              
                        ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  ��  CFourier        -./0               
         ��                   ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  ��  CACpz        	                
                       ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  ��  CDCtf         � � � � �                
                       ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  ��  CDCsens         � � � �                 
                       ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j                  ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  ��  CShow         1              
                       ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  ��  CShowmod         2              
                       ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  �� 
 CLinearize        M�  ����        ��������               
                       ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  ��  CParamTranSweep        3456789:;<=>?               
                       ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j                ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  ��  CParamACSweep        �������������               
                       ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  ��  CMonteCarlo_op        @ABCDEFGHIJKLMNOPQRSTUVWXYZ[               
                              ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  ��  CMonteCarlo_dc        \]^_`abcdefghijklmnopqrstuvw               
                       ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  ��  CMonteCarlo_ac        xyz{|}~��������������������               
                       ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  ��  CMonteCarlo_tran        ����������������������������               
                       ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  ��  CACsens        �����������               
                              ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j  ��  CNetworkAnalysis        �����������               
                       ����            P               �                        v(vout)       ����                  �                       v(4)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(2)       ����                  ء  �� �|p�|����m�|+j  ء  �� �|p�|����m�|+j                  ����            P                 >           ��   CDigSimResTemplate                ���       ����  ����:�0�yU>20.00n���   ����                       Arial����                       Arial����                       Arial  �   �  �                                ����  ���� ������       ����  ���� ������                 �               ����  �����       200������         0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial      �       �         �     �   �  �  Circuit1                  ����  ��    ��������                                                                                             �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            Z  �                5 5�� �� 5 5E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                      �  �                ��         �  @                  ���                                                  �  @  #�     <   �  <     ��                                                        #�     |   �  |     ��                                                        #�     �   �  �     ��                                                        #�     �   �  �     ��                                                        H� �      �  4     ��                                                      �      �  4   �      �  4   [title]                                       H� �   D   �  t     ��                                                      �   D   �  t   �   D   �  t   [description]                                       H� `   �   h  �     ��                                                      `   �   h  �   `   �   h  �   [id]                                       H� �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       H�      �   8    ��        	                                                   �   8       �   8  Date :         �  X  �                  H� �     �  4   	 ��        
                                              �     �  4  �     �  4  [date]                                       H�       t   8    
 ��                                                            t   8         t   8   Title :         �  0  �                  H�    L   �   x     ��                                                         L   �   x      L   �   x   Description :         �  �  X                  H�    �   �   �     ��                                                         �   �   �      �   �   �   ID :         d  �                    H�    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :         $  H  �                   ��������������          �     	title box    Analog Misc      �?    9 
 ߀     M�  ����        ��������M�  ����       ��������M�  ����       ��������M�  ����       ��������M�  ����       ��������        9                                      ������� ����     �            title                �            description               �            id               �            designer               �            date                           ����            `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                                                                                            2         �  �              � � �                   ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                          �   ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    
cgs 76         47 80moh5.6 
Q22_ 27mvrd nmodel npn_gene_g     �                      TIME� # ) time                      �                        v(3)      v(3)    TIME                 �                        v(4)      v(4)    TIME                 �                       v(vout)      v(vout)    TIME                           2         �  �           Time  � � �             np_g    ����                       Arial����                       Arial                              ����  �����z�`?2.035181e-003��G�6      ����  �����z�`?2.035181e-003��G�6      ����  ����1��{��%�-1.075922e+001������      ����  ����1��{��%�-1.075922e+001������                                                                                                                                                                                                                                                                                                                                                                                                                               1m  0                            100   100                                                             1m  0                            100   100                                1m  0                            100   100                                1m  0                            100   100                                                 
                 1m  0                            100   100                                ��   CMiniPartPin    ����11     PAS1�      �   ����22     PAS2�     BatteryBattery                          �    ����GndGnd     GNDGnd}      GndGnd                  �    ����C+C+     PASC+�      �   ����C-C-     PASC-�     capacitor_genericcapacitor_generic                          �    ����R+R+     PASR+      �   ����R-R-     PASR-     resistor_genericresistor_generic                          �    ����VCCvcc     PASVCC:      �   ����	THRESHOLDthr     PAS	THRESHOLD;     �   ����Controlctrl     PASControl<     �   ����TRIGGERtrg     PASTRIGGER=     �   ����RESETrst     PASRESET>     �   ����	DISCHARGEdis     PAS	DISCHARGE?     �   ����OUTPUTout     PASOUTPUT@     �   ����GROUNDground     PASGROUNDA     ua555ua555                                                                          �    ����MM       ��������MarkerMarker                                                                                                                                                                                                                                                                                                                    ,�e    �f � ��e                           ��e                                        ! � ��t                                                        ����       �� <                                                                               �    �Q                        6                             B 2.    224912E-003
IOUT                           @    2 2 2 2 d                                 