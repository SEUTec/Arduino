    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz    ��  CPart    �����   �  �  �����   �  �              voltage_source��  CIntPin    ��  CWire    �        �	   /   �   �      /   �   �                  Marker ��  CExtPin    ��  CVertex   �  �   ��  CSegment    �      �    �    �      @                       �    �   �                       	        `      M     @  �          VControl     ��   CPin                   ��                                                           `   M��  TLine     P       `     ��    ���                                                 ��  TPolygon     ����    ����   ��                                                         ��  TPoint    0    �����   @     � �    P    `G��0   @    �     ��  
 TTextField       �   ,     ��                                                             �   ,         �   ,   	[refname]       X  �  �  x        �   ,                Marker     Miscellaneous      �?    +   ��   CMarkerBehavior     ��  CValue             0.0      �������� M ��  	 TModelPin ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      "   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  + 1             & Analog MiscV   Generic   VControlVControl          ����               VControl  v(VControl)  N ��   CPartPin    ����MM       A ��U����RootmarkerGeneric              VControl �      �       �   �  �      �   �  �              vcswitch�    �    + �    ,    �       �   �         �   �                 1n4007- �   �     �    0     �           �   �           �   �               Gnd1 	�    �   �  �   �   �   �  �   5         4     �   �      �   �   �   �  �   �   �   �  �   ; �   �   �  �   =         <          :     9 �   �   �  �   ?          :          8     7 �   �      �   A         8          4                 `       Gnd}   �  �          gnd1     �                    ��                                                               Gnd�                   ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��    p�Z         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         C D E G   F      Ground    
Ground DINMiscellaneous      �?       ��   CGroundBehavior       Gnd ��   CBehPin     Gnd        ����Gnd����                        ��gndgnd                 K Analog Meters   Generic   gnd1gnd1          ����  gnd '�    ����GndGnd      GNDAGnd �)����SourcesGroundGeneric              0 / �   0    �           �   �          �   �              Battery�    �    �    P    �   /   �      �   /   �      �               MarkerQ 	�    �"   �  �   �   �   �  `   U         T     �   �    �  �   W         T                `      M     `  �         VSource     �                   ��                                                           `   M�    `       `     ��    ���                                                 � ����`  ����`     ��                                                         �����`    �� �    p    
 ! �   `    @��    P    p�S    � 0   P   �   t     ��                                                       0   P   �   t   0   P   �   t   	[refname]       �  p  �          �   ,    [   Y ` Z  �
  Marker     Miscellaneous      �?    +   !�     #�             0.0      �������� M %� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     P a   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  + 1             c Analog MiscV   Generic   VSourceVSource          ����               VSource  
v(VSource)  N '�    ����MM       A p�\����RootmarkerGeneric              VSource O �    P    �       _   @  �      _   @  �              Ammeter2e �   �	    �    h  	 �       _      �      _      �              capacitor_generici �   �    k �   l   �
       �   �   �      �   �   �              resistor_generic�    h   	 n 5 m 	�    �   �	  @   �   �   �	  �    �   �   �  �    �   u �
   �  �   v  	          �   �   �  �    x �   y �   �      z  	           	   u     t  	   s     r �   s �      �    �   } �          ~  	           | �
   } �   `  �    �   � �   `  �   �  	           � �   � �&   �  �    �!   � �   �  @   �  	           �  	        	        	        	   q      	  
            �   R+  	�   �   �	  �   �   � �!   �	  �   � �   �$   �  �   � �6   �   �  �   �         �     �   � �%   �  @   �                �     �   � �#      �   �   �       �   �        �     � �	   �   `  �   �        �                        
          @  R-   �	  �         RC     �                    ��                                                           @   R+�                   ��                                                          �   R-�     �   �����     ��    ���                                                 �    �   �����     ��                                                        �    �   �����     ��    ���                                                 �    x   �����     ��    (�K                                                �    x   ����l     ��                                                       �    `       X     ��    ��K                                                �     @       X     ��                                                       �    `   ����l    	 ��        	                                                �     �       �    
 ��        
                                                �     t   �   �     ��                                                           t   �   �       t   �   �   [resistance]        
  �  �  r      `   �   �   �     @   �   d     ��                                                           @   �   d       @   �   d   	[refname]        
  @  �
  �          t   $    � � � � � � � � � � � � �  �  resistor    resistor DINMiscellaneous      �?       ��  CResistorBehavior     #� ����    �חA100meg      ��������#� ���� 27     ��������#� ����       ��������#� ����       �������� R+R- J�     R+        ����R+����                        ��J�    R-      ����R-����                        �� resistor    �           � � Passive   Generic   RCRC          ����    R '�    ����R+R+      PASAR+X�U����'�   ����R-R-      PASAR-    ����Passive Generic              3 �   l   �       �   �   �      �   �   �              resistor_generic�    �
    �   �  
 �       �     �      �     �              Inductor�    h   	 � 5 � 	�            �   L+K  	�   �	            
                 �  L-L      `          L1     �                    ��                                                           @   L+�                   ��                                                          �   L-��   TArc    �       �    
                                                           �����      �   �����      �       �       �           �� �����      �    	                                                           �����      �   �����      �       �       �           �� �����   �����                                                               ����x      �   ����x      �       �       x           �� �����   �����                                                               ����`      x   ����`      x       x       `           � ����d   ����X     ��    ���                                                 � ����X   ����d     ��                                                        � ����@   ����d     ��    ���                                                 �     @       `     ��    (�K	                                                �     �       �     ��       
                                                � $   t   �   �     ��                                                       $   t   �   �   $   t   �   �   [Inductance]       l  �  l  R      \   �   |   � $   @   �   d     ��                                                       $   @   �   d   $   @   �   d   	[refname]       l     �  �          �   $    � � �   �   �   �   � � �   �   �   �   �  �  Inductor     Miscellaneous      �?    
   ��  CInductorBehavior     #� ���       �?375m      ��������#� ���� x     �������� L+L- J�     L+        ����L+����                        ��J�    L-      ����L-����                        �� Inductor  
 T           � � Passive   Generic   L1L1          ����  L '�    ����L+L+      PASAL+B 1.����'�   ����L-L-      PASAL-��X����PassiveInductorGeneric              6 �  � J�     R+        ����R+����                        ��
 6  
 � 6 � 	�    �        �   R+  	�   �       @  R-      @         RL     �                    ��                                                           @   R+�                   ��                                                          �   R-�     �   �����     ��                                                        �    �   �����     ��                                                        �    �   �����     ��                                                        �    x   �����     ��                                                        �    x   ����l     ��                                                        �    `       X     ��                                                        �     @       X     ��                                                        �    `   ����l    	 ��        	                                                �     �       �    
 ��        
                                                �     t   �   �     ��                                                           t   �   �       t   �   �   [resistance]       `  �  �  2      `   �   �   �     @   �   d     ��                                                           @   �   d       @   �   d   	[refname]       `     �  �          t   $    � � � � � � � � � � � � �  �  resistor    resistor DINMiscellaneous      �?       ��     #� �����������?0.1      ��������#� ���� 27     ��������#� ����       ��������#� ����       �������� R+R- � J�    R-      ����R-����                        �� resistor    �           � � Passive   Generic   RLRL          ����    R '�    ����R+R+      PASAR+�I�����'�   ����R-R-      PASAR-    ����Passive Generic              3 �   l   �       S   �  ,      S   �  ,              Ammeter�    �    �   �   �       _   �  �      _   �  �              
Voltmeter2�    h   	 � 5 � 	�    �    `   `   M+    	�   �*   �  �   �   � �   �  �   �    �'   `  �   �"   �   `  `   �        �     � �#   �(      �   �         �         �     �                  `   �  M-    @  �          VRL    
 �                    ��                                                               M+�                   ��                                                          �   M-�     �       �     ��    ���                                                 �             <     ��                                                        �    $      4     ��    ���                                                 �    ,      ,     ��    (�K                                                �    �      �     ��               	FIXED_ROT                                        �� 
 TRectangle     <   �   �                  ����                                             <   �   �   �    D   �   x     ��                                                         D   �   x      D   �   x   [value]       L  �  ,  B     D   �   x   � 8      �   0    	 ��        	                                               8      �   0   8      �   0   	[refname]       �    �  �  8      �   0    � � � � �           �   � 
     Voltemeter-Vert    Voltemeter-Vert_smallMiscellaneous      �?       ��   CVoltmeterBehavior     #� ����   ���"�-9.50      �������� M+M- J� 4  M+        �  M+����                        ��J� 4  M-      �  M-����                        ��	voltmeter	voltmeter   _            Analog Meters   Generic   VRLVRL          ����  IVm '�    ����M+M+      PASAM+�7      '�   ����M-M-      PASAM-�7     Analog MetersVoltmeter-verticalGeneric              7 �   �   �       �   �   �      �   �   �              resistor_generic�    h   	 5 	�    �        �   R+  	�   �       @  R-   `            RLoad     �                    ��                                                           @   R+�                   ��                                                          �   R-�     �   �����     ��    ��)                                                �    �   �����     ��    p�Z                                                �    �   �����     ��                                                       �    x   �����     ��    D�Z                                                �    x   ����l     ��    ��d                                                �    `       X     ��    |�f                                                �     @       X     ��    <�b                                                �    `   ����l    	 ��    ��)	                                                �     �       �    
 ��        
                                                �     t   �   �     ��                                                           t   �   �       t   �   �   [resistance]       �  |  `        `   �   �   �     @   �   d     ��                                                           @   �   d       @   �   d   	[refname]       �  �  �  �          t   $     �  resistor    resistor DINMiscellaneous      �?       ��     #� ����     ��@40k      ��������#� ���� 27     ��������#� ����       ��������#� ����       �������� R+R- J�     R+        ����R+����                        ��J�    R-      ����R-����                        �� resistor    �           "#Passive   Generic   RLoadRLoad          ����    R '�    ����R+R+      PASAR+    ����'�   ����R-R-      PASAR-8Lk����Passive Generic              7 �  #J� �  M+        R  M+����                        �� 7   � 7 � 	�    �    �  �   M+    	�   �       �   M-    `            V_IRL    	 �                   ��                                                       �   @   M+�                   ��                                                          @   M-�    @       @     ��    ���                                                 � �   @   �   @     ��                                                        � �   (   �   (     ��    ���                                                  � �         d                   ����                                               �   d   � �����   �����     ��          @ @                                           �|   (    
JV1��   0    G7 *��        9054@ @ � (   4   �   \     ��                                                      (   4   �   \   (   4   �   \   [value]       �  �    R  $   $   �   L   �     �����        ��                                                           �����          �����      	[refname]       �  �  �  �      �����       .  )3*  -  4/,  +	   Ammeter    Ammeter_smallMiscellaneous      �?       ��   CAmmeterBehavior     #� �i   ��tw? 5.73m      �������� M+M- &J� �  M-      R  M-����                        ��AmmeterAmmeter   _            &8Analog Meters   Generic   V_IRLV_IRL          ����  VAm '�    ����M+M+      PASAM+        '�   ����M-M-      PASAM-       Analog MetersAmmeterGeneric              3 �   l   * 3  J�    C-      ����C-����                        ��J�    2      ����2����                        ��� � 8 3   j 3 	�    �       �  C-�  	�   w        �   C+�   �            C1     �                   ��                                                           �   C-�                   ��                                                          @   C+�     @       �      ��    ���                                                 �     �   �����     ��    x�                                                 �     �   �����     ��    ���                                                 �     �       �     ��    (�K                                                � 0   t   �   �     ��                                                       0   t   �   �   0   t   �   �   [capacitance]       p  |  	        `   �   �   � 0   @   �   d     ��                                                       0   @   �   d   0   @   �   d   	[refname]       p  �  �  �          �   $    BCDEF    G      @A �  	Capacitor     Miscellaneous      �?       ��  CCapacitorBehavior     #� '  T�qs*�>24u      ��������#� ����      �?1     ��������#� ����       ��������#� ����       �������� C+C- J�     C+        ����C+����                        ��< 	capacitor   T           N<Passive   Generic   C1C1          ����  C '�    ����C+C+      PASAC+0258����'�   ����C-C-      PASAC-000E����Passive Generic              5 g o � �  N� J�    M-      ����M-����                        ��� "	 5 	 f 5 	�    X    `   �  M+2  	�   {   `   `   M-3   `  �         	V_ISource    	 �                    ��                                                           �   M+�                   ��                                                              M-�     �       �     ��                                                        �     <             ��                                                         � @   <   �����                  ����                                         ����<   @   �   � ����x   ����L     ��                                                        �  ������� �������  ��          @ @                                           �����H    ��b�����T    
>DA�����T    uT@ @ � ����D   <   |     ��                                                      ����D   <   |   ����D   <   |   [value]       4  l  �       D   �   |   �    �����        ��                                                          �����         �����      	[refname]       l  �  L  (     �����      
 TUVWX^  Y_Z	   Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       5�     #� `���   �w��-937.73n      �������� M+M- J�     M+        ����M+����                        ��QAmmeterAmmeter   V            bQAnalog Meters   Generic   	V_ISource	V_ISource          ����  VAm '�    ����M+M+      PASAM+8�W����'�   ����M-M-      PASAM-��W����Analog MetersAmmeter-verticalGeneric              VSource  J�     1       ����1����                        ��bc  VSource   N VSource M 	�    V    `       1�  	�   >   `   �  2�   `  `          X1     �                    ��                                                               1�                   ��                                                          �   2�             $     ��    ��)                                                �     \       �     ��                                                        �    8   0   8    	 ��    ��)                                                �     H   @   H     ��    p�Z                                                �     $   @   $     ��                                                       �    \   0   \     ��    D�Z                                                �               ���                                                      �               ���   �Z	                                                � `          $    
 ��        
                                               `          $   `          $   	[devname]        ����������������`          $   � `   $      H     ��                                                       `   $      H   `   $      H   	[refname]       �  �  �  l  `   $      H    hijknopq    rs    m  l     Battery     Miscellaneous      �?    9 
 ��  CParamSubBehavior     #� ����      (@12      �������� 12 eJ�    2      ����2����                        ��BatteryBattery
 9 i             ewSources   Generic   X1X1          ������   CParamSubModelType��    BATTERY2.SUBCKT Xbattery 1 2
V1 1 2 DC {voltage}
.ENDS
   ��  	 CParmDefn    1battery voltage   ParamSubvoltageV                X '�    ����11      PASA10Ab����'�   ����22      PASA2�1b����SourcesBatteryGeneric              0 �   0     0 �   0    * 0 �    0     �           �   �           �   �               Gnd�	�    �4   �  �   �'   �5   �  �   �&   �/   �  @   �        �    �     �    �(   ��6   �  �   ��)   �2   �  `   �        �                         `       Gndj   @  �          gnd2     �                    ��                                                               Gnd�                   ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��    ���          AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         ����  �     Ground    
Ground DINMiscellaneous      �?       H�       Gnd J�     Gnd        ����Gnd����                        ��gndgnd                 �Analog Meters   Generic   gnd2gnd2          ����  gnd '�    ����GndGnd      GNDAGnd�������SourcesGroundGeneric              0 �   0    �       �   @  @      �   @  @              CCVS�    �    �    �   �       �      �      �      �              Multiplier Block (XSpice)��   �    ��    �   �       �   @  @      �   @  @              VCVS��   0    �0 	�    �1   �      �   �3   �  `   ��%   ��-      `   �               �                   �  S+
G6 	�   �      �  S-URCE �  �         E2_VRL    
 �                   ��                                                           �   S+�                   ��                                                          @  S-�     �       �     ��                                                        �            @    ��                                                        �    �   �����     ���                                                       �     �       �     ���                                                       � �����      �     ��                	FIXED_ROT                                        � ����`   ����`      ��                                                         �    �        �@   �        �            ������            � P   �     �     ��                                                       P   �     �   P   �     �   	[devname]        ����������������    �����      � P   �     �    	 ��        	                                               P   �     �   P   �     �   	[refname]       �  �  0  \         �   8    �  ����    ���  �  �
 �  Controlled Voltage Source     Miscellaneous      �?       ��  CVCVSBehavior     #� ����      �?1��    ��������#� ���� VRL     �������� V+V- J� �8  V+        �  V+����                        ��J� �8  V-      �  V-����                        ��J�  �8  VC+      �   ����                        ��J�  �8  VC-      �   ����                        ��VCVSVCVS                 ����Sources   Generic   E2_VRLE2_VRL          ���� ����      �?1��    ��������VRL    E '�    ����S+V+      PASAS+        '�   ����S-V-      PASAS-P�1   SourcesVoltage Controlled Voltage SouGeneric              12  J� �7  in2����   �  in2����                        ��� 12  �12 �   �    �    �   �   /   �   �      /   �   �                  Marker�	�    �P   �      �5   �+   �      �        �    �,   �.          �       �               `      M�EX    �          PRL     �                   ��                                                           `   M�     P       `     ��                                                       �     ����    ����   ��                                                         �    0        �   @      �    P       �0   @            � ���������   !     ��                                                       ���������   !   ���������   !   	[refname]       �  �  v  w        �   ,    �  ���     Marker     Miscellaneous      �?    +   !�     #�             0.0      �������� M %� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     ��  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  + �            �Analog MiscV   Generic   PRLPRL          ����               PRL  v(PRL)  N '�    ����MM       A hQ�����RootmarkerGeneric              PRL �    �   �       �      �      �      �              Integrator Block (XSpice)��   �    �    �   �   /   �   �      /   �   �                  Marker�	�    �7   �      �*   �)   �
      �       �    �7   ��L   �  @   �   ��O      @   �            �                   `      M     @  �          Int_PRL     �                   ��                                                           `   M�     P       `     ��    ���                                                 �     ����    ����   ��                                                         �    0        �   @      �    P       �0   @            � ���������   !     ��                                                       ���������   !   ���������   !   	[refname]       �
  �  >  w        �   ,    �  ���     Marker     Miscellaneous      �?    +   !�     #�             0.0      �������� M %� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     ��  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  + �            �Analog MiscV   Generic   Int_PRLInt_PRL          ����               Int_PRL  
v(Int_PRL)  N '�    ����MM       A     ����RootmarkerGeneric              Int_PRL ��    �   �       �      @      �      @              Divider Block (XSpice)��   �    �    �   �   /   �   �      /   �   �                  Marker�	�    �@   �      �9   ��K   @      ��2   �9   �
      �       �    �:   �J   @      �8   ��N          �           �    �                       `      M     @  �          Int_PSource     �                   ��                                                           `   M�     P       `     ��                                                        �     ����    ����   ��                                                         �    0        �   @      �    P       �0   @            � ���������   !     ��                                                       ���������   !   ���������   !   	[refname]       �
  �    w        �   ,      �      Marker     Miscellaneous      �?    +   !�     #�             0.0      �������� M %� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     �  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  + �            	Analog MiscV   Generic   Int_PSourceInt_PSource          ����               Int_PSource  v(Int_PSource)  N '�    ����MM       A I QM����RootmarkerGeneric              Int_PSource �   �  �       �      �      �      �              Integrator Block (XSpice)�    �    �       �   /   �   �      /   �   �                  Marker	�    �Q   �      �4   �:   �                  �1   �<                                `      M
>DA    �          PSource     �                   ��                                                           `   M�     P       `     ��    
G6                                                 �     ����    ����   ��                                                         �    0        �   @      �    P       �0   @            � ���������   !     ��                                                       ���������   !   ���������   !   	[refname]       �  �  >  w        �   ,           Marker     Miscellaneous      �?    +   !�     #�             0.0      �������� M %� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �       �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  + �            !Analog MiscV   Generic   PSourcePSource          ����               PSource  
v(PSource)  N '�    ����MM       A  �U����RootmarkerGeneric              PSource �     �       �      �      �      �              Multiplier Block (XSpice)�    �    %�    &   �       �   @  @      �   @  @              CCVS'�   0    (0 	�    �A   �      �3   +�0          ,                           �  S+VSOU	�   �B   �  @   �    /�R   �  �   �-   1�?   �  �   2�$   3�S   �  �   �.   �>   �  `   6        5    4                      0                       �  S-7
NE �  �         H2    
 �                   ��                                                           �   S+�                   ��                                                          @  S-�     �       �     ��    ���:                                                �            @    ��    NE2_                                                �    �   �����     ���    �k                                                �     �       �     ���    �3�                                                � �����      �     ��    ���        	FIXED_ROT                                        � ����`   ����`      ��                                                         �    �        �@   �        �        SOUR������    # �     � P   �     �     ��                                                       P   �     �   P   �     �   	[devname]        ����������������    �����      � P   �     �    	 ��        	                                               P   �     �   P   �     �   	[refname]       �  �  P  <         �   8    ?  9:;>    DE=  <  8
 �  Controlled Voltage Source     Miscellaneous      �?       ��  CCCVSBehavior     #� ����      �?1��    ��������#�@ ���� 	V_ISource     �������� H+H- J� 9  H+        �  H+����                        ��J� :  H-      �  H-����                        ��CCVSCCVS                 JKRoot   Generic   H2H2          ���� ����      �?1��    ��������	V_ISource  H '�    ����S+H+      PASAS+ �     '�   ����S-H-      PASAS- �@
   SourcesCurrent Controlled Voltage SouGeneric              13  J� �7  in1����    �  in1����                        ��J 13   $13 �   �    O�    P   �       �   @  @      �   @  @              VCVSQ�   0    R0 	�    �=   �      �/   �T   �  `   �0   W�;      `   X           V    U                   �  S+��	�   7      �  S-RL.I �  �         E1    
 �                   ��                                                           �   S+�                   ��                                                          @  S-�     �       �     ��    4?
G                                                �            @    ��    
NE2                                                �    �   �����     ���   3 �                                                �     �       �     ���   I �P                                                � �����      �     ��     #O�        	FIXED_ROT                                        � ����`   ����`      ��                                                         �    �        �@   �        �            ������            � P   �     �     ��                                                       P   �     �   P   �     �   	[devname]        ����������������    �����      � P   �     �    	 ��        	                                               P   �     �   P   �     �   	[refname]       �  �  0  \         �   8    b  \]^a    gh`  _  [
 �  Controlled Voltage Source     Miscellaneous      �?       ��     #� ����      �?1��    ��������#� ���� VSource     �������� V+V- J� �8  V+        �  V+����                        ��J� �8  V-      �  V-����                        ��J�  �8  VC+      �   ����                        ��J�  �8  VC-      �   ����                        ��VCVSVCVS                 lmnoSources   Generic   E1E1          ���� ����      �?1��    ��������VSource    E '�    ����S+V+      PASAS+NDDA    '�   ����S-V-      PASAS-IRL    SourcesVoltage Controlled Voltage SouGeneric              14  J� �7  in2����   �  in2����                        ��l 14  $14 #	�    -          in1VSOU	�   Y      �  in2;
NE	�           out?
G7    �          A4     �                    ��                                                           `   in1�                   ��                                                          �   in2�                   ��                                                         `   out �     @   �   �                  ����                                             @   �   �   �     `       `     ��    5438                                                �     �       �     ��    G8 �                                                � �   `      `     ��    RL.I                                                � (   P   p   p     ��                                                      (   P   p   p   (   P   p   p   in1       �  �    R  (   P   p   p   � (   p   p   �     ��                                                      (   p   p   �   (   p   p   �   in2       �  0    �  (   p   p   �   � �   P   �   p    	 ��        	                                              �   P   �   p   �   P   �   p   out       �  �  0  R  �   P   �   p   �     �����       
 ��        
                                                   �����          �����      	[devname]        ����������������    �����      �        �   <     ��                                                              �   <          �   <   	[refname]       �  (     �         �   <    vwxyz{|}~��     Multiplier Block (XSpice)     Miscellaneous      �?    8   ��  CXSpiceBehavior       in1in2out NrJ� �7  out����   �  out����                        ��Multiplier Block (XSpice)Multiplier Block (XSpice)  8 S            Nr�Analog MiscV   Generic   A4A4                 * time value  A '�    ����in1in1      PASAin1�:
G    '�   ����in2in2      PASAin2RCE.   '�   ����outout      PASAoutG6 >   Analog Miscmultiplier blockGeneric              PSource  �J� �7  in����    �  in����                         ��! PSource   PSource 	�              in %`	�   �        outURCE �  �          A3    	 �                    ��                                                           `   in�                   ��                                                         `   out� �   `      `     ��    ~%?                                                 �     @   �   �                  ����                                             @   �   �   �     `       `     ��    �~%?                                                � (   P   p   p     ��                                                      (   P   p   p   (   P   p   p   in       X  �  �  R  (   P   p   p   � �   P   �   p     ��                                                      �   P   �   p   �   P   �   p   out       x	  �  �	  R  �   P   �   p   �     �����        ��                                                           �����          �����      	[devname]        ����������������    �����      �        �   <     ��                                                              �   <          �   <   	[refname]       @  (  �  �         �   <   	 ���������	     Integrator Block (XSpice)     Miscellaneous      �?    8   ��       inout �J� �7  out����   �  out����                        ��Integrator Block (XSpice)Integrator Block (XSpice)  8 S            ��Analog MiscV   Generic   A3A3                 * time value  A '�    ����inin      PASAin��     '�   ����outout      PASAout �    Analog Miscintegrator blockGeneric              Int_PSource � �	J� �7  den����   Z  den����                         �� Int_PSource  �Int_PSource �   �    �    �   �   /   �      �   /   �      �               Marker�	�    �I      �                   `      M	   �  �         	Rendiment     �                   ��                                                           `   M� 0   `       `     ��                                                        � ����@   ����@      ��                                                         �P   `        �@   P      �0   `       �@   p            � `   P      t     ��                                                       `   P      t   `   P      t   	[refname]       �  p  �    ���������   !    �  ��� �  Marker     Miscellaneous      �?    +   !�     #�             0.0      �������� M %� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     ��  �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  + �            �Analog MiscV   Generic   	Rendiment	Rendiment          ����               	Rendiment  v(Rendiment)  N '�    ����MM       A Pg����RootmarkerGeneric              	Rendiment � J� �7  out����   Z  out����                        ��� 	Rendiment  �	Rendiment 	�    �          num    	�   �      �  den   	�   �     �  out                  A5     �                    ��                                                           `   num�                   ��                                                          �   den�                   ��                                                         �   out �     @   �   �                  ����                                             @   �   �   �     `       `     ��    ���                                                 �     �       �     ��    t�U                                                � �   �      �     ��    ���                                                 � (   P   p   p     ��                                                      (   P   p   p   (   P   p   p   num       �    @  �  (   P   p   p   � (   �   p   �     ��                                                      (   �   p   �   (   �   p   �   den       �  �  (  R  (   �   p   �   � �   p   �   �    	 ��        	                                              �   p   �   �   �   p   �   �   out       �  p  `  �  �   p   �   �   �     �����       
 ��        
                                                   �����          �����      	[devname]        ����������������    �����      �        �   <     ��                                                              �   <          �   <   	[refname]       �  h              �   <    ������������     Divider Block     Miscellaneous      �?    8   ��       numdenout J� �7  num����    Z  num����                         ����Divider Block (XSpice)Divider Block (XSpice)  8               ���Analog MiscV   Generic   A5A5                 * time value  A '�    ����numnum      PASAnum8��    '�   ����denden      PASAden0   '�   ����outout      PASAout��>   Analog Miscdivider blockGeneric              Int_PRL  J� �7  out����   �  out����                        ���� Int_PRL  �Int_PRL 	�    �          in    	�   �        out    �  �          A1    	 �                    ��                                                           `   in�                   ��                                                         `   out� �   `      `     ��                                                        �     @   �   �                  ����                                             @   �   �   �     `       `     ��    ��K                                                � (   P   p   p     ��                                                      (   P   p   p   (   P   p   p   in       X  �  �  R  (   P   p   p   � �   P   �   p     ��                                                      �   P   �   p   �   P   �   p   out       x	  �  �	  R  �   P   �   p   �     �����        ��                                                           �����          �����      	[devname]        ����������������    �����      �        �   <     ��                                                              �   <          �   <   	[refname]       @  (  �  �         �   <   	 ���������	     Integrator Block (XSpice)     Miscellaneous      �?    8   ��       inout J� �7  in����    �  in����                         ���Integrator Block (XSpice)Integrator Block (XSpice)  8 S            ��Analog MiscV   Generic   A1A1                 * time value  A '�    ����inin      PASAin        '�   ����outout      PASAout       Analog Miscintegrator blockGeneric              PRL � �J� �7  out����   �  out����                        ��� PRL  �PRL 	�    �,          �+   �8   �      �        �                      in1    	�   �      �  in2   	�   �        out       �          A2     �                    ��                                                           `   in1�                   ��                                                          �   in2�                   ��                                                         `   out �     @   �   �                  ����                                             @   �   �   �     `       `     ��    ��K                                                �     �       �     ��    ��K                                                � �   `      `     ��    ���                                                 � (   P   p   p     ��                                                      (   P   p   p   (   P   p   p   in1       �  �    R  (   P   p   p   � (   p   p   �     ��                                                      (   p   p   �   (   p   p   �   in2       �  0    �  (   p   p   �   � �   P   �   p    	 ��        	                                              �   P   �   p   �   P   �   p   out       �  �  0  R  �   P   �   p   �     �����       
 ��        
                                                   �����          �����      	[devname]        ����������������    �����      �        �   <     ��                                                              �   <          �   <   	[refname]       �  (     �         �   <    ������������     Multiplier Block (XSpice)     Miscellaneous      �?    8   ��       in1in2out J� �7  in1����    �  in1����                        ����Multiplier Block (XSpice)Multiplier Block (XSpice)  8 S            ���Analog MiscV   Generic   A2A2                 * time value  A '�    ����in1in1      PASAin1        '�   ����in2in2      PASAin2@      '�   ����outout      PASAout       Analog Miscmultiplier blockGeneric              E_IRL � �J� 9  H+        �  H+����                        �� E_IRL   �E_IRL �	�    �       �  S+    	�   �      �  S-    �  �         H1    
 �                   ��                                                           �   S+�                   ��                                                          @  S-�     �       �     ��    ���                                                 �            @    ��                                                        �    �   �����     ���   ���                                                 �     �       �     ���   (�K                                                � �����      �     ��               	FIXED_ROT                                        � ����`   ����`      ��                                                         �    �        �@   �        �        SOUR������    # �     � P   �     �     ��                                                       P   �     �   P   �     �   	[devname]        ����������������    �����      � P   �     �    	 ��        	                                               P   �     �   P   �     �   	[refname]       �  �  P  <         �   8    �  ����    ���  �  �
 �  Controlled Voltage Source     Miscellaneous      �?       F�     #� ����      �?1��    ��������#�@ ���� V_IRL     �������� H+H- �J� :  H-      �  H-����                        ��CCVSCCVS                 ��Root   Generic   H1H1          ���� ����      �?1��    ��������V_IRL  H '�    ����S+H+      PASAS+>END    '�   ����S-H-      PASAS-�C�9   SourcesCurrent Controlled Voltage SouGeneric              0 ��    0     �           �   �           �   �               Gnd�	�    3   `       Gnd     @  �          gnd3     �                    ��                                                               Gnd�                   ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ                Ground    
Ground DINMiscellaneous      �?       H�       Gnd J�     Gnd        ����Gnd����                        ��gndgnd                 Analog Meters   Generic   gnd3gnd3          ����  gnd '�    ����GndGnd      GNDAGndJ}p�����SourcesGroundGeneric              0 )S J�    V-      ����V-����                        ��wK J�    4      ����4����                        ��J�    D-      ����D-����                        �����mK  0   . 0 	�    �   �  �                           D+   	�   6       @  D-    �  �         D1     �                   ��                                                           `   D+�                   ��                                                          �   D-�     �       �      ��    ���                                                 �     �   �����     ��                                                        �     �   �����     ��    ���                                                 �     `       �     ��                                                       �    �       �     ��    ��K                                                �     �   �����     ��    ��K                                                �     �       �     ��    N D                                                � 0   `   �   �    	 ��        	                                               0   `   �   �   0   `   �   �   	[devname]        �������������������������      � 0   �   �   �    
 ��        
                                               0   �   �   �   0   �   �   �   	[refname]       p  \  �  �  ����   �   <                   �  diode     Miscellaneous      �?       ��  CDiodeBehavior     #� ����        ��������#� ���� 27     ��������#� ����       ��������#� ����       �������� D+D- J�     D+        ����D+����                        ��d1n4007d1n4007    �          !Diode   Generic   D1D1                D '�    ����D+D+      PASAA�d?
����'�   ����D-D-      PASAK]����DiodeDiode	FairchildDO-41             8  J�     1       ����1����                        ��! 8   * 8 ;) 	�       �   �  1S  	�   �   �      2T  	�             3U  	�   B       �  4V               X2     �                    ��                                                       @   �   1�                   ��                                                      @   `   2�                   ��                                                          `   3�                   ��                                                          �   4�     �       �     ��    ��                                                �     `       �     ��                                                        �     �       �    
 ���   ��                                                � �����      �    	 ���   p�H                                                ��  TEllipse <   �   D   �                  ����                                         <   �   D   �   <   �   D   �    � �����      �               	   ����                                         �����      �   � @   `   @   �     ��       
                                                � 0   �   @   �     ��    D�H                                                � @   �   @   �     ��                                                       � �����      �     ��  � �H        	FIXED_ROT                                        �    �   4   �     ��                                                        � T   �   �   �     ��                                                       T   �   �   �   T   �   �   �   	[refname]         �  �  |      (   t   L   � �   �   4  �     ��                                                       T   `   �   �   T   `   �   �   	[devname]        ����������������       �   (    )*+,346      .7  809:5-/    2 �
  vcswitch     Miscellaneous      �?   9 
 t�    #� ����333333@4.8      ��������#� ����433333�?0.3     ��������#�  ʚ;�������?0.1     ��������#� ����    �cA10meg     �������� 1234 $=J�    3      ����3����                        ��vcswitchvcswitch
 9               $=@Switches   Generic   X2X2          ����x���voltage controlled switch   VCSW{.subckt vcsw 1 2 3 4
S 1 2 3 4 switch
.model switch sw (vt={(Von+Voff)/2} vh={(Von-Voff)/2} ron={Ron} roff={Roff})
.ends   z�    1turnon voltage   ParamSubVon               z�    1turnoff voltage   ParamSubVoffV             z�    0on resistance   ParamSubRonOhm             z�    0off resistance   ParamSubRoffOhm               X '�    ����11      PASA1Hx����'�   ����22      PASA2    ����'�   ����33      PASA3��Z����'�   ����44      PASA4OL  ����Switches Generic              VControl   J�     V+        ����V+����                        ��@&  VControl    VControl ~	�               V+g  	�   @       �  V-h   �  �         V1     �                   ��                                                           `   V+�                   ��                                                          �   V-1�     �   �����                   ����                                         �����       �   �����       �   �    �   �����     ��    ��)                                                �     �       �     ��    ��`                                                �     �       �     ��    ��)                                                �     \       �     ��    p�Z                                                � �����   
   �    
 ��               	FIXED_ROT                                        � \   `   \   `     ��                                                      \   `   \   `   \   `   \   `           �     �                   � 0   �   �   �     ��        	                                               0   �   �   �   0   �   �   �   [dc]       0  �  h  &          p   @   � 0   \   �   �    	 ��        
                                               0   \   �   �   0   \   �   �   	[refname]       0  �  �  �      ����t       O  PQSNRUVW      T    M �  Voltage Source    Voltage Source DINRoot      �?       ��  CVSourceBehavior     #� ����        0      ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       �������� V+V- J
volt_sourcevolt_source   +0            J
Sources   Generic   V1V1          ����       #�0            0      ��������#�0����      @5     ��������#�0            0     ��������#�0P�  �h㈵��>5u     ��������#�0P�  �h㈵��>5u     ��������#�0 Zb����Mbp?4m     ��������#�0 ��{�G�z�?20m     ��������    #�0            0      ��������#�0����      @5     ��������#�0����     ��@10k     ��������#�0            0     ��������#�0            0     ��������    #�0            0      ��������#�0����      �?1     ��������#�0����      �?1     ��������#�0            0     ��������#�0����      �?1     ��������    #�0            0      ��������#�0����      �?1     ��������#�0            0     ��������#�0 N  �����>2u     ��������#�0'  ���ư>1u     ��������#�0'  ���ư>1u     ��������    #�  ���� 0 0      ��������                0      �������� ����       �������� ����       �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������               V '�    ����V+V+      PWR+AV+NDDA����'�   ����V-V-      PWR-AV- � ����Sources Generic              j N � 2 � f * .  n � R � ��$����R �(���   0  P ����l h � � , ��&P; ; ; � � r 5 ��9 � 7 � � | ; v U ? z = � t �  W A x � ~ �   � � 0� � � 4��������26VX�,�� ����U N U X > @ � �  � 4 � w � 8 6 �   V B s � : <  q  � } u y { � � � T � � � � � � �� �����-���������YU73�+/            ����  ���15W   ��  CLetter    IRC modela les perdues al Condensador.
RL modela les perdues al Inductor.�	  �  �  �	     
����Arial����                       Arial     ��   �Per C=1.3u, RC=1meg, L=1.15 H i RL=0.5 ohms aquest circuit s'estabilitza als 4 o 5 segons.
Per valors m�s gras de RC S'estabilitza m�s promte.
Per RL m�s petites tamb�, s'estabilitza m�s promte.�   /
  �  �      ����Arial����                       Arial     ��   9Per RL massa petites la tensi� de sortida no �s senoidal.w     �        ����Arial����                       Arial     ��   �Amb condensadors m�s grans i inductancies m�s petites, podem incrementar la potencia.
Per� necesita m�s temps per a estabilitzarse.�    �  �      ����Arial����                       Arial            
 #�@ ����        ��������#�             0     ��������#� ����      @5     ��������#�  ʚ;�������?.1     ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true
     ��������#� ����  false     ��������               
                  #� ����        ��������#� ����       ��������#�  ����       ��������#�@ ����       ��������#�@ ����       ��������               
                  #� ����        ��������#� ����       ��������#�@ ����       ��������#�  ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������               
                 #� ����dec     ��������#� ����     @�@1k     ��������#� ����    ��.A1meg     ��������#� ����       20     ��������#� ���� true     ��������#� ���� true     ��������#� ���� true	     ��������#� ����  false
     ��������               
                 #�  ����        ��������#�  ����       ��������#�  ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������               
                  	 #� ����        ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������               
                 #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
                    #�             0      ��������#� ����      @3000m     ��������#� @KL ����Mb@?0.5m     ��������#� @KL ����Mb@?0.5m     ��������#� ���� True     ��������#� ����  F     ��������#� ���� true     ��������#� ����  false     ��������               
                 #� ����     @�@1K      ��������#�  ����       ��������#�  ����       ��������#�  ����       ��������               
         ��              #�  ����        ��������              
                  #�  ����        ��������              
                                  
                 #�  ���� RLoad      ��������#�  ���� 
resistance     ��������#� ����     @�@1k     ��������#� ����     ��@10k     ��������#� ����     @�@1k     ��������#�             0     ��������#� ����      �?500m     ��������#� @B -C��6?0.1m     ��������#� @B -C��6?0.1m     ��������#� ���� True	     ��������#� ����  false
     ��������#� ���� true     ��������#� ����  false     ��������               
                 #� ����       5      ��������#� ����       5     ��������#� ����       5     ��������#� ����       5     ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#�@ ����       ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#� ���� true     ��������#� ���� true     ��������#� ����  false     ��������#� ���� true     ��������#� ����  false      ��������#� ���� true!     ��������#� ����  false"     ��������               
                        #� ����       5      ��������#� ����       5     ��������#� ����       5     ��������#� ����       5     ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#�@ ����       ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#� ���� true     ��������#� ���� true     ��������#� ����  false     ��������#� ���� true     ��������#� ����  false      ��������#� ���� true!     ��������#� ����  false"     ��������               
                 #� ����       5      ��������#� ����       5     ��������#� ����       5     ��������#� ����       5     ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#�@ ����       ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#� ���� true     ��������#� ���� true     ��������#� ����  false     ��������#� ���� true     ��������#� ����  false      ��������#� ���� true!     ��������#� ����  false"     ��������               
                 #� ����       5      ��������#� ����       5     ��������#� ����       5     ��������#� ����       5     ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#�@ ����       ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#� ���� true     ��������#� ���� true     ��������#� ����  false     ��������#� ���� true     ��������#� ����  false      ��������#� ���� true!     ��������#� ����  false"     ��������               
                 #�@ ����        ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����decade     ��������#� ���� true     ��������#� ���� true     ��������#� ���� true     ��������#� ����  false     ��������               
                 #� ����        ��������#� ����       ��������#�@ ����       ��������#�  ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������               
                        #� ����dec     ��������#� ����     @�@1k     ��������#� ����    ��.A1meg     ��������#� ����       20     ��������#� ����        0     ��������#� ����        0     ��������#� ���� true	     ��������#� ���� true
     ��������#� ����      I@50     ��������#� ���� true     ��������#� ����  false     ��������               
                         / #� ���� x'     ��������#�     �-���q=1E-12     ��������#� @B -C��6?1E-4     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x	     ��������#� ���� x!     ��������#� ����    �  500
     ��������#� ���� x     ��������#� ����    �  500     ��������#� ���� x$     ��������#� ���� x$     ��������#� ���� x%     ��������#� ���� x"     ��������#�  ���� x*     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x&     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x+     ��������#� ���� x,     ��������#� ���� x-     ��������#� ���� xg     ��������#� ���� xf     ��������#� ���� xd     ��������#� ���� xe     ��������#� ���� xh     ��������#� ���� xj     ��������#� ���� xi     ��������#� ���� xk     ��������#� ����    e��A1Gl     ��������#�             0�     ��������#� ����      @5�     ��������#� ����      @2.5�     ��������#� ����      �?.5�     ��������#� ����      @4.5�     ��������#� 
   ��&�.>1n�     ��������#� 
   ��&�.>1n�     ��������#� 
   ��&�.>1n�     ��������#� 
   ��&�.>1n�     ��������           ��  CPrimitiveModel    d1n4007   #�    1�a��%>2.55e-9      ��������#� ���� 27     ��������#�  �/�$��?0.042     ��������#� ����      �?1.75     ��������#�  �  ��v��(�>5.76e-6     ��������#�     �]}IW�=1.85e-11     ��������#� ����      �?0.75     ��������#� ����Zd;�O�?0.333     ��������#� ���� 1.11	     ��������#� ���� 3.0
     ��������#�      0     ��������#� ���� 1     ��������#� ���� 0.5     ��������#� ����     @�@1000     ��������#� � Ǯ���?9.86e-5     ��������     Diode Generic��   CPrimitiveModelType Junction Diode model����DD   z����� 1.0E-14Saturation current    ProcessisAmp0       e     z����� 27!Parameter measurement temperature    ProcesstnomDeg C0     s     z����� 0Ohmic resistance    ProcessrsOhm0      f     z����� 1Emission Coefficient    Processn 0      g     z����� 0Transit Time    Processttsec0     h     z����� 0Junction capacitance    ProcesscjoF0     i     z����� 0     Processcj0F0     i     z����� 1Junction potential    ProcessvjV0      j     z����� 0.5Grading coefficient    Processm 0      k     z����� 1.11Activation energy    ProcessegeV0     	 l     z����� 3.0#Saturation current temperature exp.    Processxti 0     
 m     z����� 0flicker noise coefficient    Processkf 0      t     z����� 1flicker noise exponent    Processaf 0      u     z����� 0.5#Forward bias junction fit parameter    Processfc 0      n     z����� infReverse breakdown voltage    ProcessbvV0      o     z����� 1.0e-3$Current at reverse breakdown voltage    ProcessibvA0      p     z�����  Ohmic conductance    ProcesscondMho     r        D����   integrator_block2 8  #�      0.0      ��������#� ���� 1.0     ��������#� ���� -1t     ��������#� ���� 1t     ��������#� '   1u     ��������#�      0.0     ��������     integrator block Generic��2 integrator block3   INTEGRATOR_BLOCKA   z�3    0.0input offset3   Process	in_offset               z�3    1.0gain3   Processgain              z�3    -1toutput lower limit3   Processout_lower_limit             z�3    1toutput upper limit3   Processout_upper_limit             z�3    1uupp & lower sm. range3   Processlimit_range              z�3    0.0output initial condition3   Processout_ic                 int  ��   
mult_block= 8  #�      	[0.0 0.0]      ��������#�      	[1.0 1.0]     ��������#� ���� 1.0     ��������#�      0.0     ��������     multiplier block Generic��= multiplier block8   
MULT_BLOCKA   z�8    	[0.0 0.0]input offset array8   Process	in_offset              z�8    	[1.0 1.0]input gain array8   Processin_gain             z�8    1.0output gain8   Processout_gain              z�8    0.0output offset8   Process
out_offset                 mult  ��   divider_block- 8 	 #�      0.0      ��������#� ���� 1.0     ��������#�      0.0     ��������#� ���� 1.0     ��������#�     .1n     ��������#�      .1f     ��������#� ���� false     ��������#� ���� 1.0     ��������#�      0.0     ��������ӥ   divider block Generic��- divider block,   DIVIDER_BLOCKA	   z�,    0.0numerator offset,   Process
num_offset               z�,    1.0numerator gain,   Processnum_gain              z�,    0.0denominator offset,   Process
den_offset              z�,    1.0denominator gain ,   Processden_gain              z�,    .1ndenominator lower limit,   Processden_lower_limit              z�,    .1fdenominator smoothing domain,   Process
den_domain              z�,    false(smoothing fraction/absolute value switch,   Processfraction              z�,    1.0output gain,   Processout_gain              z�,    0.0output offset ,   Process
out_offset                 divide       u;                Ariald     h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j                   ����             �r               ��  TSignal                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                      v(vrl)       ����                  �                     i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CDCsweep       
 ����������               
                       ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                       v(vrl)       ����                  �                      i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACsweep        ��������               
                       ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                      v(vrl)       ����                  �                     i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  �� 
 CTranSweep       ��������               
                       ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                       v(vrl)       ����                  �                      i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACdisto        �����               
                           ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                       v(vrl)       ����                  �                      i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  9�        #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
         �                 ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                       v(vrl)       ����                  �                      i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  9�        #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
                           ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                       v(vrl)       ����                  �                      i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  9�        #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
                           ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                       v(vrl)       ����                  �                      i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  9�        #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
         �                 ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                       v(vrl)       ����                  �                      i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  9�        #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
                       	    ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                       v(vrl)       ����                  �                      i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACnoise        ��������               
                    
    ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                      v(vrl)       ����                  �                     i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  Ņ         #�  ����        ��������#�  ����       ��������#�  ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������              
                        ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                      v(vrl)       ����                  �                     i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CFourier        ����               
         ��                   ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                      v(vrl)       ����                  �                     i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACpz        	 ���������               
                       ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                      v(vrl)       ����                  �                     i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CDCtf         �����               
                       ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                      v(vrl)       ����                  �                     i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CDCsens         �����������               
                       ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                       v(vrl)       ����                  �                      i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j                  ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                      v(vrl)       ����                  �                     i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CShow         �              
                       ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                      v(vrl)       ����                  �                     i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CShowmod         �              
                       ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                      v(vrl)       ����                  �                     i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  �� 
 CLinearize        #�  ����        ��������               
                       ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                      v(vrl)       ����                  �                     i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CParamTranSweep        �������������               
                       ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                      v(vrl)       ����                  �                     i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  �              ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                       v(vrl)       ����                  �                      i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CParamACSweep        HIJKLMNOPQRST               
                       ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                      v(vrl)       ����                  �                     i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CMonteCarlo_op        ����������������������������               
                              ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                      v(vrl)       ����                  �                     i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CMonteCarlo_dc        ������������ 	
               
                       ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                       v(vrl)       ����                  �                      i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CMonteCarlo_ac         !"#$%&'()*+               
                       ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                      v(vrl)       ����                  �                     i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CMonteCarlo_tran        ,-./0123456789:;<=>?@ABCDEFG               
                       ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                       v(vrl)       ����                  �                      i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACsens        UVWXYZ[\]^_               
                              ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                       v(vrl)       ����                  �                      i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CNetworkAnalysis        `abcdefghij               
                       ����            P               �                        v(vcontrol)       ����                  �                       
v(vsource)       ����                  �                       
v(int_prl)       ����                  �                       v(int_psource)       ����                  �                       
v(psource)       ����                  �                       v(prl)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �	                       v(7)       ����                  �
                       v(8)       ����                  �                       v(e_irl)       ����                  �                       v(12)       ����                  �                       v(13)       ����                  �                       v(14)       ����                  �                       i(v1)       ����                  �                       v(vrl)       ����                  �                      i(v_isource)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j                  ����            P                 >           ��   CDigSimResTemplate                ���       ����  ����:�0�yU>20.00n���   ����                       Arial����                       Arial����                       Arial  �   �  �                                ����  ���� ������       ����  ���� ������                 �               ����  �����       200������         0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial      �       �         �     �   �  �  Circuit1                  ����  ��    ��������                                                                                                                     g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     ��   CPackageAliasSuperPCBStandardDIODE3      G�Eagle	DIODE.LBRDO41-7   AC  G�Orcad 	DAX2/DO41      G�	Ultiboard	L7DIO.l55DIO_DO41              A                                                                                                                                                                                                                                                                                                                    �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            p  �                R E� �� N AE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                      �  �                 �         �  @                  ���                                                  �  @  �     <   �  <     ��                                                        �     |   �  |     ��                                                        �     �   �  �     ��                                                        �     �   �  �     ��                                                        � �      �  4     ��                                                      �      �  4   �      �  4   [title]                                       � �   D   �  t     ��                                                      �   D   �  t   �   D   �  t   [description]                                       � `   �   h  �     ��                                                      `   �   h  �   `   �   h  �   [id]                                       � �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       �      �   8    ��        	                                                   �   8       �   8  Date :       �    H
  �                  � �     �  4   	 ��        
                                              �     �  4  �     �  4  [date]                                       �       t   8    
 ��                                                            t   8         t   8   Title :       �     
  �                  �    L   �   x     ��                                                         L   �   x      L   �   x   Description :       �  �  �  �                  �    �   �   �     ��                                                         �   �   �      �   �   �   ID :       �  �  �	  P                  �    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �  \  8                     NOPQRSTUVXYZ[\          W     	title box    Analog Misc      �?    9 
 t�     #�  ����        ��������#�  ����       ��������#�  ����       ��������#�  ����       ��������#�  ����       ��������        9                                      ����x��� ����     z�            title                z�            description               z�            id               z�            designer               z�            date                           ����            `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                                                                                            2         �  �              � � �                   ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                          �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   
cgs 76         47 80moh5.6 CE.I )Q7mvrd nmodel 
ORENDIM_P     �                       TIME� # ) time                      �                        i(v1)� < � i(v1)    TIME                 �                        v(3)      v(3)    TIME                 �                        v(5)      v(5)    TIME                 �                        v(vcontrol)      v(vcontrol)    TIME                 �                        
v(vsource)      
v(vsource)    TIME                 �    (v(5)-v(7))                  v(VRL)� �   v(VRL)    TIME                 �                        v(7)      v(7)    TIME                 �                        v(prl)      v(prl)    TIME                 �                        v(e_irl)      v(e_irl)    TIME                 �                       i(v_irl)  � � i(v_irl)    TIME                 �    i(v_irl)*v(vrl)                    PRL� � �  ����TIME                 �                        
v(int_prl)      
v(int_prl)    TIME                 �                        v(int_psource)      v(int_psource)    TIME                 �                       i(v_isource)�   � i(v_isource)    TIME                 �                        
v(psource)      
v(psource)    TIME                 �                        v(rendiment)      v(rendiment)    TIME                           2         �  �           Time  � � �           I�
H    ����                       Arial����                       Arial                              ����  ����	m9��J@2.911565e+000������      ����  ����E��S��@2.843537e+000������      ����  ������Q�^�?1.960625e+000������      ����  ����A|����-8.480212e-002��9t�                                    �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   
cgs 76                 5.6 ��������mvrd nmodel     �i��L                 2         �  �           time  � � �            E      ����                       Arial����                       Arial                              ����  ����H�]��-�?3.934240e-001������      ����  �������aeY�?3.492063e-001������      ����  �����9τ. @8.090857e+000������      ����  �����S�*���-7.710591e+000������                                                                                         �                      �                                                                                                                                                                                                                                                                                                                              �
  �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      1m  0                            100   100                                                             1m  0                            100   100                                1m  0                            100   100                                1m  0                            100   100                                                 
                 1m  0                            100   100                            ��   CPartPackage �@
 ��   CPackageg   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     HIJK      ��   CMiniPartPin    ����V+V+     PWR+V+g      ��   ����V-V-     PWR-V-h     voltage_sourcevoltage_source                          ��    ����C+C+     PASC+�      ��   ����C-C-     PASC-�     capacitor_genericcapacitor_generic                          ��    ����11     PAS1�      ��   ����22     PAS2�     BatteryBattery                          ��    ����L+L+     PASL+K      ��   ����L-L-     PASL-L     InductorInductor                          ��    ����GndGnd     GNDGnd}      GndGnd                  ��    ����M+M+     PASM+k  4  ��   ����M-M-     PASM-l  4  
Voltmeter2
Voltmeter2                          ��    ����M+M+     PASM+2      ��   ����M-M-     PASM-3     Ammeter2Ammeter2                          ��    ����11     PAS1S      ��   ����22     PAS2T     ��   ����33     PAS3U     ��   ����44     PAS4V     vcswitchvcswitch                                       } ��    ����D+D+     PASA       ��   ����D-D-     PASK       .   ��   CPackagePin 1 D+PAS  AA�� 2 D-PAS  AKDiodeDiode	Fairchild      1n4007 D1n4007D1            diode-21n40071n4007                          ��    ����MM       ��������MarkerMarker                  ��    ����R+R+     PASR+      ��   ����R-R-     PASR-     resistor_genericresistor_generic                          ��    ����R+R+     PASR+      ��   ����R-R-     PASR-     resistor_genericresistor_generic                          ��    ����MM       ��������MarkerMarker                  ��    ����R+R+     PASR+      ��   ����R-R-     PASR-     resistor_genericresistor_generic                          ��    ����M+M+     PASM+0  �  ��   ����M-M-     PASM-1  �  AmmeterAmmeter                          ��    ����inin     PASin�  �7  ��   ����outout     PASout�  �7  Integrator Block (XSpice)Integrator Block (XSpice)                          ��    ����in1in1     PASin1  �7  ��   ����in2in2     PASin2  �7  ��   ����outout     PASout  �7  Multiplier Block (XSpice)Multiplier Block (XSpice)                                  ��    ����in1in1     PASin1  �7  ��   ����in2in2     PASin2  �7  ��   ����outout     PASout  �7  Multiplier Block (XSpice)Multiplier Block (XSpice)                                  ��    ����S+V+     PASS+j  �8  ��   ����S-V-     PASS-k  �8  VCVSVCVS                          ��    ����GndGnd     GNDGnd}      GndGnd                  ��    ����MM       ��������MarkerMarker                  ��    ����inin     PASin�  �7  ��   ����outout     PASout�  �7  Integrator Block (XSpice)Integrator Block (XSpice)                          ��    ����S+H+     PASS+j  9  ��   ����S-H-     PASS-k  :  CCVSCCVS                          ��    ����S+V+     PASS+j  �8  ��   ����S-V-     PASS-k  �8  VCVSVCVS                          ��    ����GndGnd     GNDGnd}      GndGnd                  ��    ����MM       ��������MarkerMarker                  ��    ����S+H+     PASS+j  9  ��   ����S-H-     PASS-k  :  CCVSCCVS                          ��    ����MM       ��������MarkerMarker                  ��    ����MM       ��������MarkerMarker                  ��    ����numnum     PASnum  �7  ��   ����denden     PASden  �7  ��   ����outout     PASout  �7  Divider Block (XSpice)Divider Block (XSpice)                                  ��    ����MM       ��������MarkerMarker                                                                                                                                                                                                                                                            
m1     8 8 mm l=100u w                        used                                     �  � ���� �                                                                                                                                         (f    x=f � �'f                           �(f                            ,�e    �f � ��e                           ��e                                     �  � ���� �                         .I                                                                                                                                                                                                �  � ���� �                                                          >    `� ENDANAL
 DDA                        NL                             
PV    RCE.I h�7
JL1.I                         ^;                            ��
    a?
G4   �@
G3 �                          
>                            `�S    ��V�S  �V                        ��S                            �2�    �Q�R�XR��R�                        T�                            �;
    ��>
G6 �5A
MVSO                        @
NV                            ��    P   p   p   ��                           �?                             NW    � ��Ux� �                          MVSO                            ]�;
    VRL.I 1˒�
JL1.I                        I ��                            CONT      �@
>ENDDATA
>D                        V1.I                            �x�    J  \�VИPK                          P�V                              @       d   	[refname]                                                          
>    ATA
>DATAB 2.389                        PVIS                             .�     8/�     �+�                                                            _PRL    9
IPRL ��:
G8 ;                        URCE                                                                                                                                                                                            
NE2    .I O��1
JL1.I E                        ��*
                            
PVI    CE.I Hp3
LVIRL.                        ?
G7                            Z      �#T[  ���8zU                        ^                              ��Y>    ��Y>   �A^Z>   `                        ��[>                            ��3�    4�   @w^4�   @                        �5�    2 2 2 2 d                                                                                                                   