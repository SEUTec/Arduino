    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz    ��  CPart    �����   �  �  �����   �  �              voltage_source��  CIntPin    ��  CWire    �        �	   /   �   �      /   �   �                  Marker ��  CExtPin    ��  CVertex   �  �   ��  CSegment    �      �    �    �      @                       �    �   �                       	        `      M     @  �          VControl     ��   CPin                   ��                                                           `   M��  TLine     P       `     ��    ���                                                 ��  TPolygon     ����    ����   ��                                                         ��  TPoint    0    �����   @     � �    P    `G��0   @    �     ��  
 TTextField       �   ,     ��                                                             �   ,         �   ,   	[refname]       X  �  �  x        �   ,                Marker     Miscellaneous      �?    +   ��   CMarkerBehavior     ��  CValue             0.0      �������� M ��  	 TModelPin ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      "   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  + 1             & Analog MiscV   Generic   VControlVControl          ����               VControl  v(VControl)  N ��   CPartPin    ����MM       A ��U����RootmarkerGeneric              VControl �      �       �   �  �      �   �  �              vcswitch�    �    + �    ,    �       �   �         �   �                 1n4007- �   �     �    0     �           �   �           �   �               Gnd1 	�    �   �  �   �   �   �  �   5         4     �   �      �   �   �   �  �   �   �   �  �   ; �   �   �  �   =         <          :     9 �   �   �  �   ?          :          8     7 �   �      �   A         8          4                 `       Gnd}   �  �          gnd1     �                    ��                                                               Gnd�                   ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��    p�Z         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         C D E G   F      Ground    
Ground DINMiscellaneous      �?       ��   CGroundBehavior       Gnd ��   CBehPin     Gnd        ����Gnd����                        ��gndgnd                 K Analog Meters   Generic   gnd1gnd1          ����  gnd '�    ����GndGnd      GNDAGnd �)����SourcesGroundGeneric              0 / �   0    �           �   �          �   �              Battery�    �    �    P    �   /   �      �   /   �      �               MarkerQ 	�    �"   �  �   �   �   �  `   U         T     �   �    �  �   W         T                `      M     `  �         VSource     �                   ��                                                           `   M�    `       `     ��    ���                                                 � ����`  ����`     ��                                                         �����`    �� �    p    
 ! �   `    @��    P    p�S    � 0   P   �   t     ��                                                       0   P   �   t   0   P   �   t   	[refname]       �  p  �          �   ,    [   Y ` Z  �
  Marker     Miscellaneous      �?    +   !�     #�             0.0      �������� M %� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     P a   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  + 1             c Analog MiscV   Generic   VSourceVSource          ����               VSource  
v(VSource)  N '�    ����MM       A p�\����RootmarkerGeneric              VSource O �    P    �       _   @  �      _   @  �              Ammeter2e �   �    �    h   �       _      �      _      �              capacitor_generici �   �    k �   l   * 3 �   l   �
       �   �   �      �   �   �              resistor_generic�    h    o 5 n 	�    �   �	  @   �   �   �	  �    �	   �      �    �   v �   @  �    �
   x �   @  @   y             w         u �   v �          {                 t     �   �   �  �    �   ~ �
   �  �               �   �   �  �    � �   � �   �      �                ~     }     t     s     r        
            �   R+  	�   �   �	  �   �   � �!   �	  �   � �   �$   �  �   �   �   �  �   �         �     �   � �%   �  @   �            �     �     �   � �#      �   �   �       �   �        �     � �   � �   @  �   �   �   @  `   �        �     �                            
          @  R-   �	  �         RC     �                    ��                                                           @   R+�                   ��                                                          �   R-�     �   �����     ��    ���                                                 �    �   �����     ��                                                        �    �   �����     ��    ���                                                 �    x   �����     ��    (�K                                                �    x   ����l     ��                                                       �    `       X     ��    ��K                                                �     @       X     ��                                                       �    `   ����l    	 ��        	                                                �     �       �    
 ��        
                                                �     t   �   �     ��                                                           t   �   �       t   �   �   [resistance]        
  �  X  r      `   �   �   �     @   �   d     ��                                                           @   �   d       @   �   d   	[refname]        
  @  �
  �          t   $    � � � � � � � � � � � � �  �  resistor    resistor DINMiscellaneous      �?       ��  CResistorBehavior     #� ����    �cA10meg      ��������#� ���� 27     ��������#� ����       ��������#� ����       �������� R+R- J�     R+        ����R+����                        ��J�    R-      ����R-����                        �� resistor    �           � � Passive   Generic   RCRC          ����    R '�    ����R+R+      PASAR+    ����'�   ����R-R-      PASAR-X�U����Passive Generic              3 �   l   �       �   �   �      �   �   �              resistor_generic�    �    �   �   �       �     �      �     �              Inductor�    h    � 5 � 	�    |        �   L+K  	�   �	                             �  L-L      `          L1     �                    ��                                                           @   L+�                   ��                                                          �   L-��   TArc    �       �    
                                                           �����      �   �����      �       �       �           �� �����      �    	                                                           �����      �   �����      �       �       �           �� �����   �����                                                               ����x      �   ����x      �       �       x           �� �����   �����                                                               ����`      x   ����`      x       x       `           � ����d   ����X     ��    ���                                                 � ����X   ����d     ��                                                        � ����@   ����d     ��    ���                                                 �     @       `     ��    (�K	                                                �     �       �     ��       
                                                � $   t   �   �     ��                                                       $   t   �   �   $   t   �   �   [Inductance]       l  �  �  R      \   �   |   � $   @   �   d     ��                                                       $   @   �   d   $   @   �   d   	[refname]       l     �  �          �   $    � � �   �   �   �   � � �   �   �   �   �  �  Inductor     Miscellaneous      �?    
   ��  CInductorBehavior     #� ��� ffffff�?1150m      ��������#� ���� x     �������� L+L- J�     L+        ����L+����                        ��J�    L-      ����L-����                        �� Inductor  
 T           � � Passive   Generic   L1L1          ����  L '�    ����L+L+      PASAL+��X����'�   ����L-L-      PASAL-B 1.����PassiveInductorGeneric              6 �  � J�     R+        ����R+����                        �� 6   � 6 � 	�    �        �   R+  	�   �       @  R-      @         RL     �                    ��                                                           @   R+�                   ��                                                          �   R-�     �   �����     ��                                                        �    �   �����     ��                                                        �    �   �����     ��                                                        �    x   �����     ��                                                        �    x   ����l     ��                                                        �    `       X     ��                                                        �     @       X     ��                                                        �    `   ����l    	 ��        	                                                �     �       �    
 ��        
                                                �     t   �   �     ��                                                           t   �   �       t   �   �   [resistance]       `  �  �  2      `   �   �   �     @   �   d     ��                                                           @   �   d       @   �   d   	[refname]       `     �  �          t   $    � � � � � � � � � � � � �  �  resistor    resistor DINMiscellaneous      �?       ��     #� ����      $@10      ��������#� ���� 27     ��������#� ����       ��������#� ����       �������� R+R- � J�    R-      ����R-����                        �� resistor    �           � � Passive   Generic   RLRL          ����    R '�    ����R+R+      PASAR+    ����'�   ����R-R-      PASAR-�I�����Passive Generic              3 �   l   �   ����    �     ����    �                 Voltmeter2_small�    h    � 5 � 	�    z    �       M+�� 	�   �   �      M-��  �  @         VLC     �                    ��                                                       @       M+�                   ��                                                      @   `   M-� @       @         ��    ��)                                                �� 
 TRectangle �           P                  ����                                                 �   P   �    $   �   L     ��                                                         $   �   L      $   �   L   [value]       �  �  d  B  ����   |   <    � � � �     �    Voltemeter-Vert_small   	voltmeterPassive      �?       ��   CVoltmeterBehavior     #� ����   xg @ 4.25      �������� M+M- J�     M+        ����M+����                        ��J�    M-      ����M-����                        ��	voltmeter	voltmeter   _            � � Analog Meters   Generic   VLCVLC          ����  I '�    ����M+M+      PASAM+    ����'�   ����M-M-      PASAM-�)����Analog MetersVoltmeter-verticalGeneric              3  J�    C-      ����C-����                        ��� J�    2      ����2����                        ��� �  3   j 3 	�    �       �  C-�  	�   �        �   C+�   �            C1     �                   ��                                                           �   C-�                   ��                                                          @   C+�     @       �      ��    ���                                                 �     �   �����     ��    x�                                                 �     �   �����     ��    ���                                                 �     �       �     ��    (�K                                                � 0   t   �   �     ��                                                       0   t   �   �   0   t   �   �   [capacitance]       p  |  0	        `   �   �   � 0   @   �   d     ��                                                       0   @   �   d   0   @   �   d   	[refname]       p  �  �  �          �   $    � �            � �  �  	Capacitor     Miscellaneous      �?       ��  CCapacitorBehavior     #� '  kN�uϵ>1.3u      ��������#� ���� x     ��������#� ����       ��������#� ����       �������� C+C- J�     C+        ����C+����                        ���  	capacitor   T           
� Passive   Generic   C1C1          ����  C '�    ����C+C+      PASAC+000E����'�   ����C-C-      PASAC-0258����Passive Generic              5 g � � p  
� � J�    M-      ����M-����                        ���  5  f 5 	�    X    `   �  M+2  	�   �   `   `   M-3   `  �         ISource    	 �                    ��                                                           �   M+�                   ��                                                              M-�     �       �     ��                                                        �     <             ��                                                        � @   <   �����                  ����                                         ����<   @   �   � ����x   ����L     ��                                                        �  ������� �������  ��          @ @                                           �����H    ��b�����T    
>DA�����T    uT@ @ � ����D   <   |     ��                                                      ����D   <   |   ����D   <   |   [value]       4  l  D       D   �   |   �    �����        ��                                                          �����         �����      	[refname]       l  �  �  (     �����      
   	   Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       ��   CAmmeterBehavior     #� j�      V�> 6.46u      �������� M+M- J�     M+        ����M+����                        ��AmmeterAmmeter   V            Analog Meters   Generic   ISourceISource          ����  VAm '�    ����M+M+      PASAM+��W����'�   ����M-M-      PASAM-8�W����Analog MetersAmmeter-verticalGeneric              VSource  J�     1       ����1����                        ��c  VSource   N VSource M 	�    V    `       1�  	�   >   `   �  2�   `  `          X1     �                    ��                                                               1�                   ��                                                          �   2�             $     ��    ��)                                                �     \       �     ��                                                        �    8   0   8    	 ��    ��)                                                �     H   @   H     ��    p�Z                                                �     $   @   $     ��                                                       �    \   0   \     ��    D�Z                                                �               ���                                                      �               ���   �Z	                                                � `          $    
 ��        
                                               `          $   `          $   	[devname]        ����������������`          $   � `   $      H     ��                                                       `   $      H   `   $      H   	[refname]       �  �  �  l  `   $      H    %&'(+,-.    /0    *  )     Battery     Miscellaneous      �?    9 
 ��  CParamSubBehavior     #� ����      @5      �������� 12 "J�    2      ����2����                        ��BatteryBattery
 9 i             "4Sources   Generic   X1X1          ������   CParamSubModelType��    BATTERY2.SUBCKT Xbattery 1 2
V1 1 2 DC {voltage}
.ENDS
   ��  	 CParmDefn    1battery voltage   ParamSubvoltageV                X '�    ����11      PASA1�1b����'�   ����22      PASA20Ab����SourcesBatteryGeneric              0 �   0     0 �   0    * 0  J�    V-      ����V-����                        ��4K J�    4      ����4����                        ��J�    D-      ����D-����                        ��  0   . 0 	�    �   �  �                           D+   	�   6       @  D-    �  �         D1     �                   ��                                                           `   D+�                   ��                                                          �   D-�     �       �      ��    ���                                                 �     �   �����     ��                                                        �     �   �����     ��    ���                                                 �     `       �     ��                                                       �    �       �     ��    ��K                                                �     �   �����     ��    ��K                                                �     �       �     ��    N D                                                � 0   `   �   �    	 ��        	                                               0   `   �   �   0   `   �   �   	[devname]        �������������������������      � 0   �   �   �    
 ��        
                                               0   �   �   �   0   �   �   �   	[refname]       p  \  �  �  ����   �   <    EFGHIJK    LM          CD �  diode     Miscellaneous      �?       ��  CDiodeBehavior     #� ����        ��������#� ���� 27     ��������#� ����       ��������#� ����       �������� D+D- J�     D+        ����D+����                        ��?d1n4007d1n4007    �          T?Diode   Generic   D1D1                D '�    ����D+D+      PASAA]����'�   ����D-D-      PASAK�d?
����DiodeDiode	FairchildDO-41             7  J�     1       ����1����                        ��T 7   * 7 m ) <	�    A   �   �  1S  	�   �   �      2T  	�             3U  	�   B       �  4V               X2     �                    ��                                                       @   �   1�                   ��                                                      @   `   2�                   ��                                                          `   3�                   ��                                                          �   4�     �       �     ��    ��                                                �     `       �     ��                                                        �     �       �    
 ���   ��                                                � �����      �    	 ���   p�H                                                ��  TEllipse <   �   D   �                  ����                                         <   �   D   �   <   �   D   �   � �����      �               	   ����                                         �����      �   � @   `   @   �     ��       
                                                � 0   �   @   �     ��    D�H                                                � @   �   @   �     ��                                                       � �����      �     ��  � �H        	FIXED_ROT                                        �    �   4   �     ��                                                        � T   �   �   �     ��                                                       T   �   �   �   T   �   �   �   	[refname]         �  �  |      (   t   L   � �   �   4  �     ��                                                       T   `   �   �   T   `   �   �   	[devname]        ����������������       �   (    \]^_fgi      aj  kclmh`b    e �
  vcswitch     Miscellaneous      �?   9 
 1�    #� ����333333@4.8      ��������#� ����433333�?0.3     ��������#� ����      �?0.5     ��������#� ����    ��.A1meg     �������� 1234 W� J�    3      ����3����                        ��>vcswitchvcswitch
 9               W� s>Switches   Generic   X2X2          ����5���voltage controlled switch   VCSW{.subckt vcsw 1 2 3 4
S 1 2 3 4 switch
.model switch sw (vt={(Von+Voff)/2} vh={(Von-Voff)/2} ron={Ron} roff={Roff})
.ends   7�    1turnon voltage   ParamSubVon               7�    1turnoff voltage   ParamSubVoffV             7�    0on resistance   ParamSubRonOhm             7�    0off resistance   ParamSubRoffOhm               X '�    ����11      PASA1��Z����'�   ����22      PASA2@
J����'�   ����33      PASA3    ����'�   ����44      PASA4Hx����Switches Generic              VControl   J�     V+        ����V+����                        ��s&  VControl    VControl ;	�               V+g  	�   @       �  V-h   �  �         V1     �                   ��                                                           `   V+�                   ��                                                          �   V-d�     �   �����                   ����                                         �����       �   �����       �   �    �   �����     ��    ��)                                                �     �       �     ��    ��`                                                �     �       �     ��    ��)                                                �     \       �     ��    p�Z                                                � �����   
   �    
 ��               	FIXED_ROT                                        � \   `   \   `     ��                                                      \   `   \   `   \   `   \   `           �     �                   � 0   �   �   �     ��        	                                               0   �   �   �   0   �   �   �   [dc]       0  �  h  &          p   @   � 0   \   �   �    	 ��        
                                               0   \   �   �   0   \   �   �   	[refname]       0  �  �  �      ����t       �  ��������      �    � �  Voltage Source    Voltage Source DINRoot      �?       ��  CVSourceBehavior     #� ����        0      ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       �������� V+V- }=volt_sourcevolt_source   +0            }=Sources   Generic   V1V1          ����       #�0            0      ��������#�0����      @5     ��������#�0            0     ��������#�0P�  �h㈵��>5u     ��������#�0P�  �h㈵��>5u     ��������#�0��� ����MbP?1m     ��������#�0�/��q����?7.8m     ��������    #�0            0      ��������#�0����      @5     ��������#�0����     ��@10k     ��������#�0            0     ��������#�0            0     ��������    #�0            0      ��������#�0����      �?1     ��������#�0����      �?1     ��������#�0            0     ��������#�0����      �?1     ��������    #�0            0      ��������#�0����      �?1     ��������#�0            0     ��������#�0 N  �����>2u     ��������#�0'  ���ư>1u     ��������#�0'  ���ư>1u     ��������    #�  ���� 0 0      ��������                0      �������� ����       �������� ����       �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������               V '�    ����V+V+      PWR+AV+ � ����'�   ����V-V-      PWR-AV-NDDA����Sources Generic              j N � 2 � f * .  o � R    0  P l h � ,          s 5    9 � 7 u y � ;  U ? � = w } �  W A � � { � �  � � & $ & X > @ A  z  � 4 � � � 8 6    | V B t � : <  r  x v ~ � � � � � T � � �    ��  CLetter    IRC modela les perdues al Condensador.
RL modela les perdues al Inductor.O  �  (  �	     
����Arial����                       Arial     ��   �Per C=1.3u, RC=1meg, L=1.15 H i RL=0.5 ohms aquest circuit s'estabilitza als 4 o 5 segons.
Per calors m�s gras de RC S'estabilitza m�s promte.
Per RL m�s petites tamb�, s'estabilitza m�s promte.   /
    �      ����Arial����                       Arial            
 #�@ ����        ��������#�             0     ��������#� ����      @5     ��������#�  ʚ;�������?.1     ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true
     ��������#� ����  false     ��������               
                  #� ����        ��������#� ����       ��������#�  ����       ��������#�@ ����       ��������#�@ ����       ��������               
                  #� ����        ��������#� ����       ��������#�@ ����       ��������#�  ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������               
                 #� ����dec     ��������#� ����     @�@1k     ��������#� ����    ��.A1meg     ��������#� ����       20     ��������#� ���� true     ��������#� ���� true     ��������#� ���� true	     ��������#� ����  false
     ��������               
                 #�  ����        ��������#�  ����       ��������#�  ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������               
                  	 #� ����        ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������               
                 #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
                    #�             0      ��������#� ����      �?1000m     ��������#� @B -C��6?0.1m     ��������#� @B -C��6?0.1m     ��������#� ���� True     ��������#� ����  F     ��������#� ���� true     ��������#� ����  false     ��������               
                 #� ����     @�@1K      ��������#�  ����       ��������#�  ����       ��������#�  ����       ��������               
         ��              #�  ����        ��������              
                  #�  ����        ��������              
                                  
                 #�@ ����        ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true	     ��������#� ����  false
     ��������#� ���� true     ��������#� ����  false     ��������               
                 #� ����       5      ��������#� ����       5     ��������#� ����       5     ��������#� ����       5     ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#�@ ����       ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#� ���� true     ��������#� ���� true     ��������#� ����  false     ��������#� ���� true     ��������#� ����  false      ��������#� ���� true!     ��������#� ����  false"     ��������               
                        #� ����       5      ��������#� ����       5     ��������#� ����       5     ��������#� ����       5     ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#�@ ����       ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#� ���� true     ��������#� ���� true     ��������#� ����  false     ��������#� ���� true     ��������#� ����  false      ��������#� ���� true!     ��������#� ����  false"     ��������               
                 #� ����       5      ��������#� ����       5     ��������#� ����       5     ��������#� ����       5     ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#�@ ����       ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#� ���� true     ��������#� ���� true     ��������#� ����  false     ��������#� ���� true     ��������#� ����  false      ��������#� ���� true!     ��������#� ����  false"     ��������               
                 #� ����       5      ��������#� ����       5     ��������#� ����       5     ��������#� ����       5     ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#�@ ����       ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ���� true     ��������#� ���� true     ��������#� ���� true     ��������#� ����  false     ��������#� ���� true     ��������#� ����  false      ��������#� ���� true!     ��������#� ����  false"     ��������               
                 #�@ ����        ��������#�@ ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����decade     ��������#� ���� true     ��������#� ���� true     ��������#� ���� true     ��������#� ����  false     ��������               
                 #� ����        ��������#� ����       ��������#�@ ����       ��������#�  ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������#� ����       ��������               
                        #� ����dec     ��������#� ����     @�@1k     ��������#� ����    ��.A1meg     ��������#� ����       20     ��������#� ����        0     ��������#� ����        0     ��������#� ���� true	     ��������#� ���� true
     ��������#� ����      I@50     ��������#� ���� true     ��������#� ����  false     ��������               
                         / #� ���� x'     ��������#�     �-���q=1E-12     ��������#� @B -C��6?1E-4     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x	     ��������#� ���� x!     ��������#� ����    �  500
     ��������#� ���� x     ��������#� ����    �  500     ��������#� ���� x$     ��������#� ���� x$     ��������#� ���� x%     ��������#� ���� x"     ��������#�  ���� x*     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x&     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x     ��������#� ���� x+     ��������#� ���� x,     ��������#� ���� x-     ��������#� ���� xg     ��������#� ���� xf     ��������#� ���� xd     ��������#� ���� xe     ��������#� ���� xh     ��������#� ���� xj     ��������#� ���� xi     ��������#� ���� xk     ��������#� ����    e��A1Gl     ��������#�             0�     ��������#� ����      @5�     ��������#� ����      @2.5�     ��������#� ����      �?.5�     ��������#� ����      @4.5�     ��������#� 
   ��&�.>1n�     ��������#� 
   ��&�.>1n�     ��������#� 
   ��&�.>1n�     ��������#� 
   ��&�.>1n�     ��������           ��  CPrimitiveModel    d1n4007   #�    1�a��%>2.55e-9      ��������#� ���� 27     ��������#�  �/�$��?0.042     ��������#� ����      �?1.75     ��������#�  �  ��v��(�>5.76e-6     ��������#�     �]}IW�=1.85e-11     ��������#� ����      �?0.75     ��������#� ����Zd;�O�?0.333     ��������#� ���� 1.11	     ��������#� ���� 3.0
     ��������#�      0     ��������#� ���� 1     ��������#� ���� 0.5     ��������#� ����     @�@1000     ��������#� � Ǯ���?9.86e-5     ��������     Diode Generic��   CPrimitiveModelType Junction Diode model����DD   7����� 1.0E-14Saturation current    ProcessisAmp0       e     7����� 27!Parameter measurement temperature    ProcesstnomDeg C0     s     7����� 0Ohmic resistance    ProcessrsOhm0      f     7����� 1Emission Coefficient    Processn 0      g     7����� 0Transit Time    Processttsec0     h     7����� 0Junction capacitance    ProcesscjoF0     i     7����� 0     Processcj0F0     i     7����� 1Junction potential    ProcessvjV0      j     7����� 0.5Grading coefficient    Processm 0      k     7����� 1.11Activation energy    ProcessegeV0     	 l     7����� 3.0#Saturation current temperature exp.    Processxti 0     
 m     7����� 0flicker noise coefficient    Processkf 0      t     7����� 1flicker noise exponent    Processaf 0      u     7����� 0.5#Forward bias junction fit parameter    Processfc 0      n     7����� infReverse breakdown voltage    ProcessbvV0      o     7����� 1.0e-3$Current at reverse breakdown voltage    ProcessibvA0      p     7�����  Ohmic conductance    ProcesscondMho     r        D��     2n                Ariald     ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j                   ����            �@               ��  TSignal                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                      v(vlc)       ����                  �                     
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CDCsweep       
 ����������               
                       ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                       v(vlc)       ����                  �                      
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CACsweep        ��������               
                       ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                      v(vlc)       ����                  �                     
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  �� 
 CTranSweep       ��������               
                       ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                       v(vlc)       ����                  �                      
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CACdisto        �����               
                           ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                       v(vlc)       ����                  �                      
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  �        #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
                           ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                       v(vlc)       ����                  �                      
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  �        #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
                           ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                       v(vlc)       ����                  �                      
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  �        #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
                           ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                       v(vlc)       ����                  �                      
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  �        #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
                           ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                       v(vlc)       ����                  �                      
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  �        #� ����        ��������#� ����       ��������#� ����       ��������#� ����dec     ��������#� ����       ��������               
                       	    ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                      v(vlc)       ����                  �                     
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CACnoise        ��������               
                    
    ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                      v(vlc)       ����                  �                     
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  f�         #�  ����        ��������#�  ����       ��������#�  ����       ��������#� ����dec     ��������#� ����       ��������#� ����       ��������#� ����  	     ��������#� ����  
     ��������              
                        ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                      v(vlc)       ����                  �                     
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CFourier        ����               
         ��                   ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                      v(vlc)       ����                  �                     
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CACpz        	 ���������               
                       ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                      v(vlc)       ����                  �                     
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CDCtf         �����               
                       ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                      v(vlc)       ����                  �                     
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CDCsens         �����������               
                       ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                       v(vlc)       ����                  �                      
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j                  ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                      v(vlc)       ����                  �                     
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CShow         �              
                       ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                      v(vlc)       ����                  �                     
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CShowmod         �              
                       ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                      v(vlc)       ����                  �                     
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  �� 
 CLinearize        #�  ����        ��������               
                       ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                      v(vlc)       ����                  �                     
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CParamTranSweep        ����                
                       ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                      v(vlc)       ����                  �                     
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  �              ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                       v(vlc)       ����                  �                      
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CParamACSweep        yz{|}~������               
                       ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                      v(vlc)       ����                  �                     
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CMonteCarlo_op        	
 !"#$               
                              ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                      v(vlc)       ����                  �                     
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CMonteCarlo_dc        %&'()*+,-./0123456789:;<=>?@               
                       ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                       v(vlc)       ����                  �                      
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CMonteCarlo_ac        ABCDEFGHIJKLMNOPQRSTUVWXYZ[\               
                       ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                      v(vlc)       ����                  �                     
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CMonteCarlo_tran        ]^_`abcdefghijklmnopqrstuvwx               
                       ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                       v(vlc)       ����                  �                      
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CACsens        �����������               
                              ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                       v(vlc)       ����                  �                      
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CNetworkAnalysis        �����������               
                       ����            P               �                        v(vcontrol)       ����                  �                       v(3)       ����                  �                       v(5)       ����                  �                       v(4)       ����                  �                       v(6)       ����                  �                       i(v1)       ����                  �                       v(vlc)       ����                  �                      
i(isource)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j                  ����            P                 >           ��   CDigSimResTemplate                ���       ����  ����:�0�yU>20.00n���   ����                       Arial����                       Arial����                       Arial  �   �  �                                ����  ���� ������       ����  ���� ������                 �               ����  �����       200������         0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial      �       �         �     �   �  �  Circuit1                  ����  ��    ��������                                                                                                                     g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     ��   CPackageAliasSuperPCBStandardDIODE3      *�Eagle	DIODE.LBRDO41-7   AC  *�Orcad 	DAX2/DO41      *�	Ultiboard	L7DIO.l55DIO_DO41              A                                                        �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            T  �                T C�� �� _ RE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                      �  �                �         �  @                  ���                                                  �  @  �     <   �  <     ��                                                        �     |   �  |     ��                                                        �     �   �  �     ��                                                        �     �   �  �     ��                                                        � �      �  4     ��                                                      �      �  4   �      �  4   [title]                                       � �   D   �  t     ��                                                      �   D   �  t   �   D   �  t   [description]                                       � `   �   h  �     ��                                                      `   �   h  �   `   �   h  �   [id]                                       � �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       �      �   8    ��        	                                                   �   8       �   8  Date :       �    H
  �                  � �     �  4   	 ��        
                                              �     �  4  �     �  4  [date]                                       �       t   8    
 ��                                                            t   8         t   8   Title :       �     
  �                  �    L   �   x     ��                                                         L   �   x      L   �   x   Description :       �  �  �  �                  �    �   �   �     ��                                                         �   �   �      �   �   �   ID :       �  �  �	  P                  �    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �  \  8                     123456789;<=>?          :     	title box    Analog Misc      �?    9 
 1�     #�  ����        ��������#�  ����       ��������#�  ����       ��������#�  ����       ��������#�  ����       ��������        9                                      ����5��� ����     7�            title                7�            description               7�            id               7�            designer               7�            date                           ����            `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                                                                                            2         �  �              � � �                   ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                          �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   
cgs 76         47 80moh5.6      
PVmvrd nmodel �
JL1.I8    	 �                      TIME� # ) time                      �                        i(v1)� < � i(v1)    TIME                 �                        v(3)      v(3)    TIME                 �    (v(5)-v(3))                  v(VLC)� �   v(VLC)    TIME                 �                        v(5)      v(5)    TIME                 �                       v(vcontrol)      v(vcontrol)    TIME                 �                        
v(vsource)      
v(vsource)    TIME                 �                      
i(isource)�   � 
i(isource)    TIME                 �    i(isource)*v(vsource)                    Pin  � �  ����TIME                           2         �  �           Time  � � �            %a    ����                       Arial����                       Arial                              ����  ����.��S��?5.804843e-001������      ����  �������z�?5.773939e-001������      ����  ������o1�i�?9.816843e-001������      ����  ���� �#G:��-5.238315e-001������                                                                         �                      �                                                                                                                                                                                                                                                                                                  �
  �
                                                                                                                                                                                                                                                                  1m  0                            100   100                                                             1m  0                            100   100                                1m  0                            100   100                                1m  0                            100   100                                                 
                 1m  0                            100   100                            ��   CPartPackage �@
 ��   CPackageg   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     +,-.      ��   CMiniPartPin    ����V+V+     PWR+V+g      [�   ����V-V-     PWR-V-h     voltage_sourcevoltage_source                          [�    ����C+C+     PASC+�      [�   ����C-C-     PASC-�     capacitor_genericcapacitor_generic                          [�    ����11     PAS1�      [�   ����22     PAS2�     BatteryBattery                          [�    ����L+L+     PASL+K      [�   ����L-L-     PASL-L     InductorInductor                          [�    ����GndGnd     GNDGnd}      GndGnd                  [�    ����M+M+     PASM+��     [�   ����M-M-     PASM-��    Voltmeter2_smallVoltmeter2_small                          [�    ����M+M+     PASM+2      [�   ����M-M-     PASM-3     Ammeter2Ammeter2                          [�    ����11     PAS1S      [�   ����22     PAS2T     [�   ����33     PAS3U     [�   ����44     PAS4V     vcswitchvcswitch                                       X [�    ����D+D+     PASA       [�   ����D-D-     PASK       .   ��   CPackagePin 1 D+PAS  AAo� 2 D-PAS  AKDiodeDiode	Fairchild      1n4007 D1n4007D1            diode-21n40071n4007                          [�    ����MM       ��������MarkerMarker                  [�    ����R+R+     PASR+      [�   ����R-R-     PASR-     resistor_genericresistor_generic                          [�    ����R+R+     PASR+      [�   ����R-R-     PASR-     resistor_genericresistor_generic                          [�    ����MM       ��������MarkerMarker                                                                                                                                                                                               
m1     8 8 mm l=100u w                        used                                     �  � ���� �                                                                                                                                         (f    x=f � �'f                           �(f                            ,�e    �f � ��e                           ��e                                     �  � ���� �                         .I                                                                                                                                                                                                �  � ���� �                                                          >    `� ENDANAL
 DDA                        NL                             
PV    RCE.I h�7
JL1.I                         ^;                            ��
    a?
G4   �@
G3 �                          
>                            `�S    ��V�S  �V                        ��S    2 2 2 2 d                                                   