    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz    ��  CPart    �����   �  �  �����   �  �              voltage_source��  CIntPin    ��  CWire    �        �   /   �   �      /   �   �                  Marker ��  CExtPin    ��  CVertex(   �  @   ��  CSegment    �   �  @                �    �+   �  �                            `      M��6               VControl     ��   CPin                   ��                                                           `   M��  TLine     P       `     ��                                                        ��  TPolygon ����   ����      ��                                                         ��  TPoint    0    �� �   @    
 ! �    P    @��0   @    p�S    ��  
 TTextField       �   ,     ��                                                             �   ,         �   ,   	[refname]       8  8  �  �        �   ,               Marker     Miscellaneous      �?    +   ��   CMarkerBehavior     ��  CValue             0.0      �������� M ��  	 TModelPin ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �          �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  + 1             $ Analog MiscV   Generic   VControlVControl          ����               VControl  v(VControl)  N ��   CPartPin    ����MM       A     ����RootmarkerGeneric              VControl �       �       �   P  @      �   P  @              irf840�    �    ) �   *    �       _      �      _      �              capacitor_generic�    �    �    .    �   ����    �     ����    �                 Voltmeter2_small/ �   *   0 3 	�    �   �  �   �   �0   �  �   4 �   �/   �
  �   �   7 �   �
  �   8             6 �   �-   �  �   �   ; �   �      <    	         : �
   �.   �  �   �   ? �   �  �   @            �   �"   �  �   B �   C �$   �  `   D                ?     >     ;         7         5         3                �       M+�� 	�   �   �  �   �	   G �!   �      H �   I �%   �
      J �   �)   �      �   �'   �  �   N    	    M     �   �   �      �   �*   �  �   R         Q     P        M     L     K     �   �,   �
  �   T         K                              �      M-��  �  �         VLC     �                    ��                                                       @       M+�                   ��                                                      @   `   M-� @       @         ��    ��)                                                �� 
 TRectangle �           P                  ����                                                 �   P   �    $   �   L     ��                                                         $   �   L      $   �   L   [value]       �    T  �  ����   |   <    V W Z [     X    Voltemeter-Vert_small   	voltmeterPassive      �?       ��   CVoltmeterBehavior     !� ����    ���?954.19m      �������� M+M- ��   CBehPin     M+        ����M+����                        ��_�    M-      ����M-����                        ��	voltmeter	voltmeter   _            ` a Analog Meters   Generic   VLCVLC          ����  I %�    ����M+M+      PASAM+�)����%�   ����M-M-      PASAM-    ����Analog MetersVoltmeter-verticalGeneric              5 �    .    �       �     �      �     �              Inductord �   �    f �    g    �
       �   �   �      �   �   �              resistor_generich �   �    j �   k   �       _   @  �      _   @  �              Ammeter2�    *    m 3 l 	�    U    `   �  M+.I �	�   �#   �
  @       
          `   `   M-V1.I �
  �         IL    	 �                    ��                                                           �   M+�                   ��                                                              M-�     �       �     ��                                                        �     <             ��                                                        Y� @   <   �����                  ����                                         ����<   @   �   � ����x   ����L     ��                                                        �  ������� �������  ��          @ @                                           �����H    ��b�����T    
>DA�����T    uT@ @ � ����D   <   |     ��                                                      ����D   <   |   ����D   <   |   [value]       T	  �  �
  B     D   �   |   � ��������b   !     ��                                                       ��������b   !   ��������b   !   	[refname]       f	  �  �	  w     �����      
 r s t u v |   w } x 	   Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       ��   CAmmeterBehavior     !� ����    ���?463.60m      �������� M+M- _�     M+        ����M+����                        ��_�    M-      ����M-����                        ��AmmeterAmmeter   V            � � Analog Meters   Generic   ILIL          ����  VAm %�    ����M+M+      PASAM+�;Q����%�   ����M-M-      PASAM-hX����Analog MetersAmmeter-verticalGeneric              7  _�    R-      ����R-����                        ���  7  i 7 	�    �   �
  �           
            �   R+  	�   q       @  R-   �
            RL     �                    ��                                                           @   R+�                   ��                                                          �   R-�     �   �����     ��    c�
                                                �    �   �����     ��     7.1                                                �    �   �����     ��    .106                                                �    x   �����     ��    0634                                                �    x   ����l     ��    O�>
                                                �    `       X     ��    G6                                                  �     @       X     ��     ��                                                �    `   ����l    	 ��    v��
	                                                �     �       �    
 ��    214E
                                                �     t   �   �     ��                                                           t   �   �       t   �   �   [resistance]       @  \  �  �      `   �   �   �     @   �   d     ��                                                           @   �   d       @   �   d   	[refname]       @  �  �  `          t   $    � � � � � � � � � � � � �  �  resistor    resistor DINMiscellaneous      �?       ��  CResistorBehavior     !� �����������?0.1      ��������!� ���� 27     ��������!� ����       ��������!� ����       �������� R+R- _�     R+        ����R+����                        ���  resistor    �           � � Passive   Generic   RLRL          ����    R %�    ����R+R+      PASAR+p����%�   ����R-R-      PASAR-�}X����Passive Generic              6  _�    L-      ����L-����                        ���  6  e 6 	�    9        �   L+K  	�   �       �  L-L   �
            L     �                    ��                                                           @   L+�                   ��                                                          �   L-��   TArc �����      �    
                                                           �����      �   �����      �       �       �           �� �����      �    	                                                           �����      �   �����      �       �       �           �� ����x      �                                                               ����x      �   ����x      �       �       x           �� ����`      x                                                               ����`      x   ����`      x       x       `           � ����d   ����X     ��    7.00                                                � ����X   ����d     ��    0016                                                � ����@   ����d     ��    2043                                                �     @       `     ��    5177	                                                �     �       �     ��    E   
                                                � $   t   �   �     ��                                                       $   t   �   �   $   t   �   �   [Inductance]       L  |  d        \   �   |   � $   @   �   d     ��                                                       $   @   �   d   $   @   �   d   	[refname]       L  �  �  �          �   $    � � �   �   �   �   � � �   �   �   �   �  �  Inductor     Miscellaneous      �?    
   ��  CInductorBehavior     !� ��� �����W?1.45m      ��������!� ���� x     �������� L+L- _�     L+        ����L+����                        ���  Inductor  
 T           � � Passive   Generic   LL          ����  L %�    ����L+L+      PASAL+�� ����%�   ����L-L-      PASAL-0HT����PassiveInductorGeneric              5 �    .    �	       �   �   �      �   �   �              resistor_generic� �   *   � 3 	�    =        �   R+  	�   O       @  R-   �  @         RC     �                    ��                                                           @   R+�                   ��                                                          �   R-�     �   �����     ��    ATA
                                                �    �   �����     ��    A
>D                                                �    �   �����     ��    >DAT                                                �    x   �����     ��    ATAB                                                �    x   ����l     ��    �W;
                                                �    `       X     ��    ;
G7                                                �     @       X     ��    G7 �                                                �    `   ����l    	 ��     ���	                                                �     �       �    
 ��    ��>

                                                �     t   �   �     ��                                                           t   �   �       t   �   �   [resistance]        	  �  8
  2      `   �   �   �     @   �   d     ��                                                           @   �   d       @   �   d   	[refname]        	     �	  �          t   $    � � � � � � � � � � � � �  �  resistor    resistor DINMiscellaneous      �?       ��     !� ����    �cA10meg      ��������!� ���� 27     ��������!� ����       ��������!� ����       �������� R+R- _�     R+        ����R+����                        ��_�    R-      ����R-����                        �� resistor    �           � � Passive   Generic   RCRC          ����    R %�    ����R+R+      PASAR+ � ����%�   ����R-R-      PASAR-�� ����Passive Generic              5 - �   .   �       _   @  �      _   @  �              Ammeter2�    �    �    �    �   /   �      �   /   �      �               Marker� 	�    �   �  `   �   �   �  �   �         �     �   � �   �  �   �                        `      M��F @  @         VSource     �                   ��                                                           `   M�    `       `     ��    ��)                                                � ����`  ����`     ��                                                         �����`    �� �    p    
 ! �   `    @��    P    p�S    � 0   P   �   t     ��                                                       0   P   �   t   0   P   �   t   	[refname]       �  0  `  �        �   ,    �   � � �  �
  Marker     Miscellaneous      �?    +   �     !�             0.0      �������� M #� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  + 1             � Analog MiscV   Generic   VSourceVSource          ����               VSource  
v(VSource)  N %�    ����MM       A  � ����RootmarkerGeneric              VSource � �    �    �           �   �          �   �              Battery� �   �     �    �     �           �   �           �   �               Gnd� 	�    �   �   
   �   �   �   
   �   �1   �   
   �   �   �   	   �         �     �      �     �          �     �   �&   �  �	   �         �                 `       Gnd}   `   
          gnd1     �                    ��                                                               Gnd�                   ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��    p�Z         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         � � � �   �      Ground    
Ground DINMiscellaneous      �?       ��   CGroundBehavior       Gnd _�     Gnd        ����Gnd����                        ��gndgnd                 Analog Meters   Generic   gnd1gnd1          ����  gnd %�    ����GndGnd      GNDAGnd �)����SourcesGroundGeneric              0 �   �     0 � �   �    �       �   �         �   �                 1n4007�    �    �     ( 4  _�    3      ����source����                        ��_�     D+        ����D+����                        �� 4   4 	�    �   �  �                          D+   	�   �       @  D-    �  �         D1     �                   ��                                                           `   D+�                   ��                                                          �   D-�     �       �      ��    ���                                                 �     �   �����     ��                                                        �     �   �����     ��    ���                                                 �     `       �     ��                                                       �    �       �     ��    ��K                                                �     �   �����     ��    ��K                                                �     �       �     ��                                                        � 0   `   �   �    	 ��        	                                               0   `   �   �   0   `   �   �   	[devname]        �������������������������      � 0   �   �   �    
 ��        
                                               0   �   �   �   0   �   �   �   	[refname]       P  <	  �  �	  ����   �   <                   �  diode     Miscellaneous      �?       ��  CDiodeBehavior     !� ����        ��������!� ���� 27     ��������!� ����       ��������!� ����       �������� D+D- 
_�    D-      ����D-����                        ��d1n4007d1n4007             
Diode   Generic   D1D1                D %�    ����D+D+      PASAA�}W����%�   ����D-D-      PASAK0vW����DiodeDiode	FairchildDO-41             0  _�    V-      ����V-����                        ��_�    2      ����2����                        ��  0   � 0 	�    �    `       1�  	�   �   `   �  2�   @  �          X1     �                    ��                                                               1�                   ��                                                          �   2�             $     ��    ��)                                                �     \       �     ��                                                        �    8   0   8    	 ��    ��)                                                �     H   @   H     ��    p�Z                                                �     $   @   $     ��                                                       �    \   0   \     ��    D�Z                                                �               ���                                                      �               ���   �Z	                                                � `          $    
 ��        
                                               `          $   `          $   	[devname]        ����������������`          $   � `   $      H     ��                                                       `   $      H   `   $      H   	[refname]       `  �  �  �  `   $      H    &'(),-./    01    +  *     Battery     Miscellaneous      �?    9 
 ��  CParamSubBehavior     !� ����      @5      �������� 12 _�     1       ����1����                        ��#BatteryBattery  9 i             5#Sources   Generic   X1X1          ������   CParamSubModelType��    BATTERY2.SUBCKT Xbattery 1 2
V1 1 2 DC {voltage}
.ENDS
   ��  	 CParmDefn    1battery voltage   ParamSubvoltageV                X %�    ����11      PASA10Ab����%�   ����22      PASA2�1b����SourcesBatteryGeneric              VSource  5� _�     M+        ����M+����                        �� VSource   � VSource � 	�    �    `   �  M+2  	�   E   `   `   M-3   @            ISource    	 �                    ��                                                           �   M+�                   ��                                                              M-�     �       �     ��                                                        �     <             ��                                                        Y� @   <   �����                  ����                                         ����<   @   �   � ����x   ����L     ��                                                        �  ������� �������  ��          @ @                                           �����H    ��b�����T    
>DA�����T    uT@ @ � ����D   <   |     ��                                                      ����D   <   |   ����D   <   |   [value]         �  �  b     D   �   |   �    �����        ��                                                          �����         �����      	[refname]       L  �  �  �     �����      
 ?@ABCI  DJE	   Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       ~�     !� bx�    +4M�-891.23u      �������� M+M- <_�    M-      ����M-����                        ��AmmeterAmmeter   V            <MAnalog Meters   Generic   ISourceISource          ����  VAm %�    ����M+M+      PASAM+8�W����%�   ����M-M-      PASAM-��W����Analog MetersAmmeter-verticalGeneric              5  ` M_�     C+        ����C+����                        ��� �  5  , 5 + 	�    S       �  C-�  	�   A        �   C+�   �  �         C     �                   ��                                                           �   C-�                   ��                                                          @   C+�     @       �      ��    282E                                                �     �   �����     ��    1E-0                                                �     �   �����     ��    -001                                                �     �       �     ��    01
J                                                � 0   t   �   �     ��                                                       0   t   �   �   0   t   �   �   [capacitance]       P  <  0  �      `   �   �   � 0   @   �   d     ��                                                       0   @   �   d   0   @   �   d   	[refname]       P  �  �  @          �   $    UVWXY    Z      ST �  	Capacitor     Miscellaneous      �?       ��  CCapacitorBehavior     !� '  H�����z>100n      ��������!� ���� x     ��������!� ����       ��������!� ����       �������� C+C- P_�    C-      ����C-����                        �� 	capacitor   T           PaPassive   Generic   CC          ����  C %�    ����C+C+      PASAC+I   ����%�   ����C-C-      PASAC-   @����Passive Generic              3 � 1 n  _�     1       ����drain����                        ��a a� �  3  ( 3 ' 	�           �  Gatew  	�   Q       �   Drainx  	�        @  Sourcey   �  `          X2     �                    ��                                                           �   Gate�                   ��                                                      `   @   Drain�                   ��                                                      `   �   Source� p   p   h   t     ��    ��)                                                � X   t   P   x     ��                                                       � X   t   h   t     ��    ��)                                                � `   @   `   �     ��    p�Z                                                � @   �   @   �     ��                                                       � ,   �   @   �     ��    �Z                                                ��  TEllipse    P   p   �    	           	                                                   P   p   �      P   p   �   � ,   \   ,   l    
 ��       
                                                � ,   x   ,   �     ��                                                        � ,   �   `   �     ��                                                        � ,   d   `   d     ��                                                        � ,   �   ,   �     ��                                                        �     `       �     ��                                                        �     �       �     ��                                                        � ����������������  ��                                                        �,   �    8�`�8   |        �8   �            � ����������������  ��                                                        �`   t    (�d�X   �    �@
>�h   �     7     � ����   �   8     ��                                                       ����   �   8   ����   �   8   	[refname]       �  �    <  ����   �   8   � ���������        ��                                                       ���������      ���������      	[devname]        �������������������������       hijklmnoprstuvwxyz~�  �     MOS 3 nmos diode     Miscellaneous      �?   #    X %�    ����Drain1      PASAD   ����%�   ����Gate2      PASAG��X����%�   ����Source3      PASASPfc����%�   ����Drain1      PASAD    ����MOSFETsPower N-channel MosfetInternational RectifierTO-220             VControl   _�     V+        ����V+����                        ��_�    2      ����gate����                        ��$  VControl    VControl 	�               V+g  	�   �       �  V-h   �  �         V1     �                   ��                                                           `   V+�                   ��                                                          �   V-q�     �   �����                   ����                                         �����       �   �����       �   �    �   �����     ��    ��)                                                �     �       �     ��    ��`                                                �     �       �     ��    ��)                                                �     \       �     ��    p�Z                                                � �����   
   �    
 ��               	FIXED_ROT                                        � \   `   \   `     ��                                                      \   `   \   `   \   `   \   `           �  �  �  �                � 0   �   �   �     ��        	                                               0   �   �   �   0   �   �   �   [dc]         0	  H  �	          p   @   � 0   \   �   �    	 ��        
                                               0   \   �   �   0   \   �   �   	[refname]         �  �  4	      ����t       �  ��������      �    � �  Voltage Source    Voltage Source DINRoot      �?       ��  CVSourceBehavior     !� ����        0      ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       �������� V+V- �"volt_sourcevolt_source   +0            �"Sources   Generic   V1V1          ����       !�0            0      ��������!�0����      @5     ��������!�0            0     ��������!�0�  I�����z>0.1u     ��������!�0�  I�����z>0.1u     ��������!�0�I iUMu�>15u     ��������!�0� :�`���?79u     ��������    !�0            0      ��������!�0����      @5     ��������!�0����     ��@10k     ��������!�0            0     ��������!�0            0     ��������    !�0            0      ��������!�0����      �?1     ��������!�0����      �?1     ��������!�0            0     ��������!�0����      �?1     ��������    !�0            0      ��������!�0����      �?1     ��������!�0            0     ��������!�0 N  �����>2u     ��������!�0'  ���ư>1u     ��������!�0'  ���ư>1u     ��������    !�  ���� 0 0      ��������                0      �������� ����       �������� ����       �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������               V %�    ����V+V+      PWR+AV+NDDA����%�   ����V-V-      PWR-AV- � ����Sources Generic              ( � � � 0 � , e � i  m    � �  * . g k                      D H > B : 6 T J  L N � �  < 8 @ � P 4 R � � � 2   2   � � Q      �       G �       �     3   � A 9 � =             I C q E K � O  M S  U ; ? 7 5 �              
 !�@ ����        ��������!�             0     ��������!� ����      @5     ��������!�  ʚ;�������?.1     ��������!�@ ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ���� true
     ��������!� ����  false     ��������               
                  !� ����        ��������!� ����       ��������!�  ����       ��������!�@ ����       ��������!�@ ����       ��������               
                  !� ����        ��������!� ����       ��������!�@ ����       ��������!�  ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������               
                 !� ����dec     ��������!� ����     @�@1k     ��������!� ����    ��.A1meg     ��������!� ����       20     ��������!� ���� true     ��������!� ���� true     ��������!� ���� true	     ��������!� ����  false
     ��������               
                 !�  ����        ��������!�  ����       ��������!�  ����       ��������!� ����dec     ��������!� ����       ��������!� ����       ��������!� ����  	     ��������!� ����  
     ��������               
                  	 !� ����        ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������               
                 !� ����        ��������!� ����       ��������!� ����       ��������!� ����dec     ��������!� ����       ��������               
                    !�             0      ��������!�  ��{�G�z�?10m     ��������!� �  I�����z>0.1u     ��������!� �  I�����z>0.1u     ��������!� ���� True     ��������!� ����  F     ��������!� ���� true     ��������!� ����  false     ��������               
                 !� ����     @�@1K      ��������!�  ����       ��������!�  ����       ��������!�  ����       ��������               
         ��              !�  ����        ��������              
                  !�  ����        ��������              
                                  
                 !�@ ����        ��������!�@ ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ���� true	     ��������!� ����  false
     ��������!� ���� true     ��������!� ����  false     ��������               
                 !� ����       5      ��������!� ����       5     ��������!� ����       5     ��������!� ����       5     ��������!� ����       ��������!� ����  	     ��������!� ����  
     ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ���� true     ��������!�@ ����       ��������!�@ ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����dec     ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ���� true     ��������!� ���� true     ��������!� ���� true     ��������!� ����  false     ��������!� ���� true     ��������!� ����  false      ��������!� ���� true!     ��������!� ����  false"     ��������               
                        !� ����       5      ��������!� ����       5     ��������!� ����       5     ��������!� ����       5     ��������!� ����       ��������!� ����  	     ��������!� ����  
     ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ���� true     ��������!�@ ����       ��������!�@ ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����dec     ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ���� true     ��������!� ���� true     ��������!� ���� true     ��������!� ����  false     ��������!� ���� true     ��������!� ����  false      ��������!� ���� true!     ��������!� ����  false"     ��������               
                 !� ����       5      ��������!� ����       5     ��������!� ����       5     ��������!� ����       5     ��������!� ����       ��������!� ����  	     ��������!� ����  
     ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ���� true     ��������!�@ ����       ��������!�@ ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����dec     ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ���� true     ��������!� ���� true     ��������!� ���� true     ��������!� ����  false     ��������!� ���� true     ��������!� ����  false      ��������!� ���� true!     ��������!� ����  false"     ��������               
                 !� ����       5      ��������!� ����       5     ��������!� ����       5     ��������!� ����       5     ��������!� ����       ��������!� ����  	     ��������!� ����  
     ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ���� true     ��������!�@ ����       ��������!�@ ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����dec     ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ���� true     ��������!� ���� true     ��������!� ���� true     ��������!� ����  false     ��������!� ���� true     ��������!� ����  false      ��������!� ���� true!     ��������!� ����  false"     ��������               
                 !�@ ����        ��������!�@ ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����decade     ��������!� ���� true     ��������!� ���� true     ��������!� ���� true     ��������!� ����  false     ��������               
                 !� ����        ��������!� ����       ��������!�@ ����       ��������!�  ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������!� ����       ��������               
                        !� ����dec     ��������!� ����     @�@1k     ��������!� ����    ��.A1meg     ��������!� ����       20     ��������!� ����        0     ��������!� ����        0     ��������!� ���� true	     ��������!� ���� true
     ��������!� ����      I@50     ��������!� ���� true     ��������!� ����  false     ��������               
                         / !� ���� x'     ��������!�     �-���q=1E-12     ��������!� @B -C��6?1E-4     ��������!� ���� x     ��������!� ���� x     ��������!� ���� x     ��������!� ���� x     ��������!� ���� x     ��������!� ���� x     ��������!� ���� x	     ��������!� ���� x!     ��������!� ����    �  500
     ��������!� ���� x     ��������!� ����    �  500     ��������!� ���� x$     ��������!� ���� x$     ��������!� ���� x%     ��������!� ���� x"     ��������!�  ���� x*     ��������!� ���� x     ��������!� ���� x     ��������!� ���� x     ��������!� ���� x&     ��������!� ���� x     ��������!� ���� x     ��������!� ���� x     ��������!� ���� x+     ��������!� ���� x,     ��������!� ���� x-     ��������!� ���� xg     ��������!� ���� xf     ��������!� ���� xd     ��������!� ���� xe     ��������!� ���� xh     ��������!� ���� xj     ��������!� ���� xi     ��������!� ���� xk     ��������!� ����    e��A1Gl     ��������!�             0�     ��������!� ����      @5�     ��������!� ����      @2.5�     ��������!� ����      �?.5�     ��������!� ����      @4.5�     ��������!� 
   ��&�.>1n�     ��������!� 
   ��&�.>1n�     ��������!� 
   ��&�.>1n�     ��������!� 
   ��&�.>1n�     ��������           ��  CPrimitiveModel    d1n4007   !�    1�a��%>2.55e-9      ��������!� ���� 27     ��������!�  �/�$��?0.042     ��������!� ����      �?1.75     ��������!�  �  ��v��(�>5.76e-6     ��������!�     �]}IW�=1.85e-11     ��������!� ����      �?0.75     ��������!� ����Zd;�O�?0.333     ��������!� ���� 1.11	     ��������!� ���� 3.0
     ��������!�      0     ��������!� ���� 1     ��������!� ���� 0.5     ��������!� ����     @�@1000     ��������!� � Ǯ���?9.86e-5     ��������     Diode Generic��   CPrimitiveModelType Junction Diode model����DD   8����� 1.0E-14Saturation current    ProcessisAmp0       e     8����� 27!Parameter measurement temperature    ProcesstnomDeg C0     s     8����� 0Ohmic resistance    ProcessrsOhm0      f     8����� 1Emission Coefficient    Processn 0      g     8����� 0Transit Time    Processttsec0     h     8����� 0Junction capacitance    ProcesscjoF0     i     8����� 0     Processcj0F0     i     8����� 1Junction potential    ProcessvjV0      j     8����� 0.5Grading coefficient    Processm 0      k     8����� 1.11Activation energy    ProcessegeV0     	 l     8����� 3.0#Saturation current temperature exp.    Processxti 0     
 m     8����� 0flicker noise coefficient    Processkf 0      t     8����� 1flicker noise exponent    Processaf 0      u     8����� 0.5#Forward bias junction fit parameter    Processfc 0      n     8����� infReverse breakdown voltage    ProcessbvV0      o     8����� 1.0e-3$Current at reverse breakdown voltage    ProcessibvA0      p     8�����  Ohmic conductance    ProcesscondMho     r        D��     3��  CMacroBehavior      123 d�	irf840irf840 #               d�	MOSFETs   International Rectifier   X2X2          ��.subckt irf840 1  2  3
**************************************
*      model generated by modpex     *
*copyright(c) symmetry design systems*
*         all rights reserved        *
*    unpublished licensed software   *
*   contains proprietary information *
*      which is the property of      *
*     symmetry or its licensors      *
*commercial use or resale restricted *
*   by symmetry license agreement    *
**************************************
* model generated on apr 29, 96
* model format: spice3
* symmetry power mos model (version 1.0)
* external node designations
* node 1 -> drain
* node 2 -> gate
* node 3 -> source
m1 9 7 8 8 mm l=100u w=100u
* default values used in mm:
* the voltage-dependent capacitances are
* not included. other default values are:
*   rs=0 rd=0 ld=0 cbd=0 cbs=0 cgbo=0
.model mm nmos level=1 is=1e-32 vto=3.84925 lambda=0.00279225 kp=6.49028 cgso=1.18936e-05 cgdo=1e-11
rs 8 3 0.0178672
d1 3 1 md
.model md d is=6.51041e-09 rs=0.0106265 n=1.49911 bv=500 ibv=0.00025 eg=1.2 xti=3.02565 tt=0.0001 cjo=1.08072e-09 vj=3.67483 m=0.9 fc=0.5
rds 3 1 2e+07
rd 9 1 0.810848
rg 2 7 3.45326
d2 4 5 md1
* default values used in md1:
*   rs=0 eg=1.11 xti=3.0 tt=0
*   bv=infinite ibv=1ma
.model md1 d is=1e-32 n=50 cjo=1.81945e-09 vj=1.07167 m=0.9 fc=1e-08
d3 0 5 md2
* default values used in md2:
*   eg=1.11 xti=3.0 tt=0 cjo=0
*   bv=infinite ibv=1ma
.model md2 d is=1e-10 n=1 rs=3e-06
rl 5 10 1
fi2 7 9 vfi2 -1
vfi2 4 0 0
ev16 10 0 9 7 1
cap 11 10 1.81945e-09
fi1 7 9 vfi1 -1
vfi1 11 6 0
rcap 6 10 1
d4 0 6 md3
* default values used in md3:
*   eg=1.11 xti=3.0 tt=0 cjo=0
*   rs=0 bv=infinite ibv=1ma
.model md3 d is=1e-10 n=1
.ends
                 Ariald        �� �|p�|����m�|+j     �� �|p�|����m�|+j                   ����            ��d              	 ��  TSignal                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                      v(vlc)       ����                  ��                     
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  ��  CDCsweep       
 ����������               
                       ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                       v(vlc)       ����                  ��                      
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  ��  CACsweep        ��������               
                       ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                      v(vlc)       ����                  ��                     
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  �� 
 CTranSweep       ��������               
                       ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                       v(vlc)       ����                  ��                      
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  ��  CACdisto        �����               
                           ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                       v(vlc)       ����                  ��                      
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  %�        !� ����        ��������!� ����       ��������!� ����       ��������!� ����dec     ��������!� ����       ��������               
                           ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                       v(vlc)       ����                  ��                      
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  %�        !� ����        ��������!� ����       ��������!� ����       ��������!� ����dec     ��������!� ����       ��������               
                           ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                       v(vlc)       ����                  ��                      
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  %�        !� ����        ��������!� ����       ��������!� ����       ��������!� ����dec     ��������!� ����       ��������               
                           ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                       v(vlc)       ����                  ��                      
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  %�        !� ����        ��������!� ����       ��������!� ����       ��������!� ����dec     ��������!� ����       ��������               
                           ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                       v(vlc)       ����                  ��                      
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  %�        !� ����        ��������!� ����       ��������!� ����       ��������!� ����dec     ��������!� ����       ��������               
                       	    ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                      v(vlc)       ����                  ��                     
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  ��  CACnoise        ��������               
                    
    ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                      v(vlc)       ����                  ��                     
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  {�         !�  ����        ��������!�  ����       ��������!�  ����       ��������!� ����dec     ��������!� ����       ��������!� ����       ��������!� ����  	     ��������!� ����  
     ��������              
                        ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                      v(vlc)       ����                  ��                     
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  ��  CFourier        �                
         ��                   ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                      v(vlc)       ����                  ��                     
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  ��  CACpz        	 ���������               
                       ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                      v(vlc)       ����                  ��                     
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  ��  CDCtf         �����               
                       ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                      v(vlc)       ����                  ��                     
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  ��  CDCsens         �����������               
                       ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                       v(vlc)       ����                  ��                      
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j                  ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                      v(vlc)       ����                  ��                     
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  ��  CShow                       
                       ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                      v(vlc)       ����                  ��                     
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  ��  CShowmod                       
                       ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                      v(vlc)       ����                  ��                     
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  �� 
 CLinearize        !�  ����        ��������               
                       ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                      v(vlc)       ����                  ��                     
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  ��  CParamTranSweep        	
               
                       ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                      v(vlc)       ����                  ��                     
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j                ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                       v(vlc)       ����                  ��                      
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  ��  CParamACSweep        �������������               
                       ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                      v(vlc)       ����                  ��                     
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  ��  CMonteCarlo_op         !"#$%&'()*+,-               
                              ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                      v(vlc)       ����                  ��                     
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  ��  CMonteCarlo_dc        ./0123456789:;<=>?@ABCDEFGHI               
                       ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                       v(vlc)       ����                  ��                      
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  ��  CMonteCarlo_ac        JKLMNOPQRSTUVWXYZ[\]^_`abcde               
                       ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                      v(vlc)       ����                  ��                     
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  ��  CMonteCarlo_tran        fghijklmnopqrstuvwxyz{|}~��               
                       ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                       v(vlc)       ����                  ��                      
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  ��  CACsens        �����������               
                              ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                       v(vlc)       ����                  ��                      
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j  ��  CNetworkAnalysis        �����������               
                       ����            P              	 ��                        
v(vsource)       ����                  ��                       v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       i(v1)       ����                  ��                       v(vlc)       ����                  ��                      
i(isource)       ����                     �� �|p�|����m�|+j     �� �|p�|����m�|+j                  ����            P                 >           ��   CDigSimResTemplate                ���       ����  ����:�0�yU>20.00n���   ����                       Arial����                       Arial����                       Arial  �   �  �                                ����  ���� ������       ����  ���� ������                 �               ����  �����       200������         0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial      �       �         �     �   �  �  Circuit1                  ����  ��    ��������                 Q   TO-220�3-Pin TO220 Package                                                                                                                                                                                                                                       �     ��   CPackageAliasSuperPCBStandardTO220      R�Orcad TO220AB      R�	UltiboardUltilib.l55TO220      R�Eagletransistor-npn.lbrTO220     R�Eagletransistor-powerTO220BV   GDS  R�Eagletransistor-powerTO220AH   BCE  R�EaglediodeTO220AB   A1A2C          A                                                                                                                                              g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     R�SuperPCBStandardDIODE3      R�Eagle	DIODE.LBRDO41-7   AC  R�Orcad 	DAX2/DO41      R�	Ultiboard	L7DIO.l55DIO_DO41              A                  �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TD                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                      �	                  Y�         �  @                  ���                                                  �  @  �     <   �  <     ��                                                        �     |   �  |     ��                                                        �     �   �  �     ��                                                        �     �   �  �     ��                                                        � �      �  4     ��                                                      �      �  4   �      �  4   [title]                                       � �   D   �  t     ��                                                      �   D   �  t   �   D   �  t   [description]                                       � `   �   h  �     ��                                                      `   �   h  �   `   �   h  �   [id]                                       � �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       �      �   8    ��        	                                                   �   8       �   8  Date :       �	  ,    �                  � �     �  4   	 ��        
                                              �     �  4  �     �  4  [date]                                       �       t   8    
 ��                                                            t   8         t   8   Title :       �	  ,  �
  �                  �    L   �   x     ��                                                         L   �   x      L   �   x   Description :       �	  �  �  �                  �    �   �   �     ��                                                         �   �   �      �   �   �   ID :       �	  �  x
  `                  �    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �	  l                         `abcdefghjklmn          i     	title box    Analog Misc      �?    9 
 2�     !�  ����        ��������!�  ����       ��������!�  ����       ��������!�  ����       ��������!�  ����       ��������        9                                      ����6��� ����     8�            title                8�            description               8�            id               8�            designer               8�            date                           ����            `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                                                                                            2         �  �              � � �                   ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                          �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   
cgs 76         47 80moh5.6 RCE.I ��mvrd nmodel �>
IL.I 91    	 ��                      TIME� # ) time                      ��                        i(v1)� < � i(v1)    TIME                 ��                        v(3)      v(3)    TIME                 ��                        
v(vsource)      
v(vsource)    TIME                 ��    (v(5)-v(3))                  v(VLC)� �   v(VLC)    TIME                 ��                        v(5)      v(5)    TIME                 ��                        v(vcontrol)      v(vcontrol)    TIME                 ��                       
i(isource)�   � 
i(isource)    TIME                 ��                      i(il)  � � i(il)    TIME                           2         �  �           Time  � � �           �t3B    ����                       Arial����                       Arial                              ����  ���� �il�?9.483564e-003����      ����  �����@`���?9.132321e-003��G{q      ����  ��������^q�?6.075892e-001������      ����  �����$f,�-5.679198e-001������                                                                         �                      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  1m  0                            100   100                                                             1m  0                            100   100                                1m  0                            100   100                                1m  0                            100   100                                                 
                 1m  0                            100   100                            ��   CPartPackage�^n	 ��   CPackageQ   TO-220�3-Pin TO220 Package                                                                                                                                                                                                                                       �     STUVWXY   ��  � ��g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     Z[\]      ��   CMiniPartPin    ����V+V+     PWR+V+g      ��   ����V-V-     PWR-V-h     voltage_sourcevoltage_source                       � ��    ����Drain1     PASDx      ��   ����Gate2     PASGw     ��   ����Source3     PASSy     ��   ����Drain1     PASDx  �   (   ��   CPackagePin 2 DrainPAS  AD�� 1 GatePAS  AG�� 3 SourcePAS  AS�� 4 DrainPAS  ADPower N-channel MosfetMOSFETsInternational Rectifier        Xirf840X1            to-220irf840irf840                                  ��    ����11     PAS1�      ��   ����22     PAS2�     BatteryBattery                          ��    ����MM       ��������MarkerMarker                  ��    ����GndGnd     GNDGnd}      GndGnd                  ��    ����M+M+     PASM+��     ��   ����M-M-     PASM-��    Voltmeter2_smallVoltmeter2_small                          ��    ����M+M+     PASM+2      ��   ����M-M-     PASM-3     Ammeter2Ammeter2                          ��    ����C+C+     PASC+�      ��   ����C-C-     PASC-�     capacitor_genericcapacitor_generic                          ��    ����L+L+     PASL+K      ��   ����L-L-     PASL-L     InductorInductor                          ��    ����R+R+     PASR+      ��   ����R-R-     PASR-     resistor_genericresistor_generic                          ��    ����R+R+     PASR+      ��   ����R-R-     PASR-     resistor_genericresistor_generic                          ��    ����MM       ��������MarkerMarker               � ��    ����D+D+     PASA       ��   ����D-D-     PASK         �� 1 D+PAS  AA�� 2 D-PAS  AKDiodeDiode	Fairchild      1n4007 D1n4007D1            diode-21n40071n4007                          ��    ����M+M+     PASM+2      ��   ����M-M-     PASM-3     Ammeter2Ammeter2                                                                                                                                                                       
m1     8 8 mm l=100u w                        used                                                                                                                                                                                            H	    �/�XF  �T                        @1                            ,�e    �f � ��e                           ��e                                     �  � ���� �                         .I                                                                                                       SOUR     ���3
JL1.I sd(<                        E                               ATA
    AB 6.9521000000E                        E.I                             <
G7    >
G6 l�@
MVSOUR                        NVCO                            L1.I    ;
G7 ����
G6 X�                        G5                              �!U    X�F�"UF  �3.                        `'U                            (f    x=f � �'f                           �(f                            5535    -004
JV1.I �	�
                        �ʽ
    2 2 2 2 d                                                     