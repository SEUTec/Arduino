    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz      ��  CPart       _   �         _   �                 capacitor_generic��  CIntPin    ��  CWire     �      �       �   �  �       �   �  �               R�    �    	 �    
    �       �   �        �   �                Inductor �   �	     �       	 �       S   �  ,      S   �  ,              Ammeter �   �    �        12  �        �   ����  �  �  ����  �  �              switch_time �   �    �      �       _   @  �      _   @  �              Ammeter2�    �     �         �           �   �           �   �               Gnd ��  CExtPin    ��  CVertex+   `  `   ��  CSegment<    �   `  `	   #         !     "�+    �J      `   % "�,    �      �   '         &          !     "�/   !  �D   �  `   "�     �K      `   "�    �6      @   -          ,     +      *     ) "�    �3   �  @   /          *                          `       Gnd}      `          gnd1     ��   CPin                    ��                                                               Gnd��  TLine                   ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        3�         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        3�    ,   4   ,     ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        3�    8   (   8     ��    p�Z         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         2 4 5 7   6      Ground    
Ground DINMiscellaneous      �?       ��   CGroundBehavior       Gnd ��   CBehPin     Gnd        ����Gnd����                        ��gndgnd                 ; Analog Meters   Generic   gnd1gnd1          ����  gnd ��   CPartPin    ����GndGnd      GNDAGnd �)����SourcesGroundGeneric              0 �       �           �   �          �   �              Battery�    �    @ �    A    �       _   @  �      _   @  �              Ammeter2B �   �    D �    E    �       _   �  �      _   �  �              
Voltmeter2F �       G 0 �     �(          "�2    �H      �   K "�5   L  �A   `  �   "�-   N  �   `  �   O            M "�4   N  �M   �  �   "�#   R  �:   �  @   S             Q "�*   R  �I      �   "�   V  �=      @   W             U                             J                `   `   M+k  �   (   `   �  M-l   �   �          IV_Vx1    
 1�                    ��                                                               M+1�                   ��                                                          �   M-3�     �       �     ��    ��                                                3�             <     ��    
NVA                                                3�    $      4     ��    ��                                                3�    ,      ,     ��    p�H                                                3�    �      �     ��               	FIXED_ROT                                        �� 
 TRectangle     <   �   �                  ����                                             <   �   �   ��  
 TTextField    D   �   x     ��                                                         D   �   x      D   �   x   [value]       �   l  �  �     D   �   x   c� 8      �   0    	 ��        	                                               8      �   0   8      �   0   	[refname]       h  �  �  o  8      �   0    Z [ ^ _ ` b d     e       ]   \ 
     Voltemeter-Vert    Voltemeter-Vert_smallMiscellaneous      �?       ��   CVoltmeterBehavior     ��  CValue ����      (@12.00      �������� M+M- :�     M+        ����M+����                        ��:�    M-      ����M-����                        ��	voltmeter	voltmeter   k            j k Analog Meters   Generic   IV_Vx1IV_Vx1          ����  IVm <�    ����M+M+      PASAM+@������<�   ����M-M-      PASAM-�����Analog MetersVoltmeter-verticalGeneric              9 �    E    �       _   @  �      _   @  �              Ammeter2n �   �    �    q    �   ����  �  �  ����  �  �              switch_timer �      s 3 �     �#   �  �   "�    �7   �  �   w        v                    �  SW+=  �    �>   �      "�(   z  �P   �  �   "�8   |  �   �  �   }             { "�$   |  �G   �  @   "�0    �Q   �  �	   "�:   �  �      �	   �            "�!   �  �F   �  �
   �            �     �      "�"   �  �8   @  @   �                                            SW->   �            X1    
 1�                   ��                                                           �   SW+1�                    ��                                                             SW-��   TArc �����                                                                      ����|       �   ����|       �       �       �           3�     �       �     ��    ���                                                 3�     �       �     ��                                                        3�     �            ��    ���                                                 3� (   �       �     ��    (�K                                                3�     �      �     ��                                                       c� 8   �   �   �     ��                                                       8   �   �   �   8   �   �   �   	[refname]       H    �  �         t   @   c� 8   |   �   �    	 ��        	                                               8   |   �   �   8   |   �   �   	[devname]        ����������������    �����       �   � � � � �   � � �   � 
 �  Switch_Open     Miscellaneous      �?   9 
 ��  CParamSubBehavior    h� ��� ����MbP?1m      ��������h� ���{�G�zt?5m     ��������h� ����      �?0.5     ��������h� ����    ��.A1meg     �������� 45 :�     4       ����4����                        ��:�    5      ����5����                        ��switch_timeswitch_time
 9               � � Switches   Generic   X1X1          ������   CParamSubModelType��time controlled switch   TIME_SWITCH�.subckt tswitch 4 5
S 4  5  3 0 switch
V0 3  0 DC 0 PWL ( 0 0
+ {time_on-.000000001} 0
+ {time_on+.000000001}  1
+ {time_off-.000000001} 1
+ {time_off+.000000001} 0)

IVm0 3  0 0

.model switch SW  vt = .5   vh = 0   ron = {res_on}   roff = {res_off}  
.ends   ��  	 CParmDefn     time the switch closes   ParamSubtime_ons              ��    1time the switch opens   ParamSubtime_offs             ��    1resistance when switch closed   ParamSubres_onOhm             ��    1megresistance when switch open   ParamSubres_offOhm               X <�    ����SW+4      PASASW+    ����<�   ����SW-5      PASASW-    ����SwitchesTime Controlled SwitchGeneric              10 p  � :�    M-      ����M-����                        �� 10  o 10 �    T    `   `   M+2  �   x   `   �  M-3   @  �          VA_X1    	 1�                    ��                                                               M+1�                   ��                                                          �   M-3�             <     ��    x�R                                                3�     �       �     ��     zT                                                a�     <   �   �                  ����                                             <   �   �   3� �   H   �   t     ��    (�K                                                ��  TPolygon ����������������  ��          @ @                                           ��  TPoint�   x    h�P���   l    �  ���   l        @ @ c�    D   �   |     ��                                                         D   �   |      D   �   |   [value]       L  �  1  :     D   �   |   c� D   ����       ��                                                       D   ����     D   ����     	[refname]         �  A  j     �����      
 � � � � � �   � � � 	     Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       ��   CAmmeterBehavior     h� n�     �|G�> 6.03u      �������� M+M- :�     M+        ����M+����                        ��� AmmeterAmmeter   �            � � Analog Meters   Generic   VA_X1VA_X1          ����  VAm <�    ����M+M+      PASAM+PǕ����<�   ����M-M-      PASAM-�������Analog MetersAmmeter-verticalGeneric              9 �    E    �       _   @  �      _   @  �              Ammeter2� �   �
    �   �  
 �       �   �         �   �                 1n4007�        � 12 � �     �9      �   "�6   �  �C      �   "�    �-   �
  �   �        �     � "�1   �  �E      @   "�%    �%    
  @   �         �     "�3   �  �O      �	   "�)    �   �  �	   �        �     � "�.   �  �N      �
   �                     �                                @  D+   �    �?      �   "�    �;      �   �  
      �      
               D-       `         D1     1�                   ��                                                           �   D+1�                   ��                                                          `   D-3� �����       �      ��    ���                                                 3�     �       �     ��                                                        3� �����       �     ��    ���                                                 3�     �       �     ��    (�K                                                3� �����       �     ��                                                       3�     �      �     ��    ��K                                                3�     �       `     ��    ��K                                                c� d   �   $  �    	 ��        	                                               0   `   �   �   0   `   �   �   	[devname]        �������������������������      c� 0   �   �   �    
 ��        
                                               0   �   �   �   0   �   �   �   	[refname]       �    9  �  ����   �   <    � � � � � � �     � �           � �  �
  diode     Miscellaneous      �?       ��  CDiodeBehavior     h� ����  F      ��������h� ���� x     ��������h� ���� x     ��������h� ���� x     �������� D+D- :�     D+        ����D+����                        ��:�    D-      ����D-����                        ��d1n4007d1n4007    �          � � Diode   Generic   D1D1                D <�    ����D+D+      PASAA   `����<�   ����D-D-      PASAK��P����DiodeDiode	FairchildDO-41             14 �  � :�    M-      ����M-����                        ��
 14 
 � 14 �    X    `   `   M+2  �   �   `   �  M-3   �  �          VA_D1    	 1�                    ��                                                               M+1�                   ��                                                          �   M-3�             <     ��    ���                                                 3�     �       �     ��                                                        a�     <   �   �                  ����                                             <   �   �   3� �   H   �   t     ��    ���                                                 �� ����������������  ��          @ @                                           ���   x    h�P���   l    �  ���   l        @ @ c�    D   �   |     ��                                                         D   �   |      D   �   |   [value]       �  �    :     D   �   |   c� D   ����       ��                                                       D   ����     D   ����     	[refname]       �  �  �  j     �����      
 � � � � � �   � � � 	     Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       ��     h� x���   ೥��-10.08m      �������� M+M- :�     M+        ����M+����                        ��� AmmeterAmmeter   �            � � Analog Meters   Generic   VA_D1VA_D1          ����  VAm <�    ����M+M+      PASAM+    ����<�   ����M-M-      PASAM-    ����Analog MetersAmmeter-verticalGeneric              9  :�    M-      ����M-����                        ��j � �  9  C 9 �     �   `  @   "�7    �   `  �                          `   �  M+2  �   P   `   `   M-3      `         VA_Ix1    	 1�                    ��                                                           �   M+1�                   ��                                                              M-3�     �       �     ��                                                        3�     <             ��                                                        a� @   <   �����                  ����                                         ����<   @   �   3� ����x   ����L     ��                                                        ��  ������� �������  ��          @ @                                           ������H    ��b������T    
>DA������T    uT@ @ c� ����D   <   |     ��                                                      ����D   <   |   ����D   <   |   [value]       �  ,  	  �     D   �   |   c� ��������O        ��                                                       ��������O      ��������O      	[refname]       �  ?    �     �����      
 	
  	   Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       ��     h� d���   @����-10.08m      �������� M+M- :�     M+        ����M+����                        �� AmmeterAmmeter   V             Analog Meters   Generic   VA_Ix1VA_Ix1          ����  VAm <�    ����M+M+      PASAM+��W����<�   ����M-M-      PASAM-8�W����Analog MetersAmmeter-verticalGeneric              4  :�     1       ����1����                        �� 4   ? 4 > �       `       1�  �   $   `   �  2�      �          XSource     1�                    ��                                                               11�                   ��                                                          �   23�             $     ��    ��)                                                3�     \       �     ��                                                        3�    8   0   8    	 ��    ��)                                                3�     H   @   H     ��    p�Z                                                3�     $   @   $     ��                                                       3�    \   0   \     ��    D�Z                                                3�               ���                                                      3�               ���   �Z	                                                c� `          $    
 ��        
                                               `          $   `          $   	[devname]        ����������������`          $   c� :   �����   ����  ��                                                       :   �����   ����:   �����   ����	[refname]       �  \  3    `   $      H     !"#    $%           Battery     Miscellaneous      �?    9 
 ��     h� ����      (@12      �������� 12 :�    2      ����2����                        ��BatteryBattery
 9 i             (Sources   Generic   XSourceXSource          ��������    BATTERY2.SUBCKT Xbattery 1 2
V1 1 2 DC {voltage}
.ENDS
   ��    1battery voltage   ParamSubvoltageV                X <�    ����11      PASA1�1b����<�   ����22      PASA20Ab����SourcesBatteryGeneric              0 H  �         �       _   @  �      _   @  �              Ammeter2-�   �    /�    0   �       �   �         �   �                 1n40071�      23 �     �L   �      "�'   5 �4   �  �   6                          @  D+   �   �          D-    �  �	         D2     1�                   ��                                                           �   D+1�                   ��                                                          `   D-3� �����       �      ��    ���                                                 3�     �       �     ��                                                        3� �����       �     ��    ���                                                 3�     �       �     ��                                                       3� �����       �     ��    ��K                                                3�     �      �     ��    ��K                                                3�     �       `     ��                                                        c� d   �   $  �    	 ��        	                                               0   `   �   �   0   `   �   �   	[devname]        �������������������������      c� 0   �   �   �    
 ��        
                                               0   �   �   �   0   �   �   �   	[refname]       0  |  �  '  ����   �   <    ;<=>?@A    BC          9: �
  diode     Miscellaneous      �?       �     h� ����  F      ��������h� ���� x     ��������h� ���� x     ��������h� ���� x     �������� D+D- :�     D+        ����D+����                        ��:�    D-      ����D-����                        ��d1n4007d1n4007    @          IJDiode   Generic   D2D2                D <�    ����D+D+      PASAA    ����<�   ����D-D-      PASAK    ����DiodeDiode	FairchildDO-41             7  :�    M-      ����M-����                        ��I 7  .7 �    0    `   �  M+2  �   7  `   `   M-3   @  `         VA_D2    	 1�                    ��                                                           �   M+1�                   ��                                                              M-3�     �       �     ��    ���                                                 3�     <             ��                                                        a�     �   �   <                  ����                                             <   �   �   3� �   x   �   L     ��    ���                                                 �� ����������������  ��          @ @                                           ���   H      � ���   T    �������   T        @ @ c�    D   �   |     ��                                                         D   �   |      D   �   |   [value]       L  ,  ^  �     D   �   |   c� E   ����       ��                                                       E   ����     E   ����     	[refname]         H  Z  �     �����      
 PQRSTZ  U[V	     Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       ��     h� X   ����?10.08m      �������� M+M- :�     M+        ����M+����                        ��MAmmeterAmmeter   �            ^MAnalog Meters   Generic   VA_D2VA_D2          ����  VAm <�    ����M+M+      PASAM+�  ����<�   ����M-M-      PASAM-���W����Analog MetersAmmeter-verticalGeneric              0  (; ^:�     M+        ����M+����                        ��k   0     0  �    .    `   �  M+2  �    �5      �   "�&    �<          e       d             `   `   M-3   �  `         VA_X2    	 1�                    ��                                                           �   M+1�                   ��                                                              M-3�     �       �     ��    ���                                                 3�     <             ��    ��K                                                a�     �   �   <                  ����                                             <   �   �   3� �   x   �   L     ��    ���                                                 �� ����������������  ��          @ @                                           ���   H      
 ���   T      ���   T        @ @ c�    D   �   |     ��                                                         D   �   |      D   �   |   [value]       �  ,  �  �     D   �   |   c� P   ����       ��                                                       P   ����     P   ����     	[refname]       �  Q  �  �     �����      
 ghijkq  lrm	     Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       ��     h� 6��    xپ-5.99u      �������� M+M- a:�    M-      ����M-����                        ��AmmeterAmmeter   �            auAnalog Meters   Generic   VA_X2VA_X2          ����  VAm <�    ����M+M+      PASAM+e"  ����<�   ����M-M-      PASAM-    ����Analog MetersAmmeter-verticalGeneric              8   u:�    5      ����5����                        �� 8   8 �    �        �  SW+=  �   f         SW->       	         X2    
 1�                   ��                                                           �   SW+1�                    ��                                                             SW-�� �����                                                                      ����|       �   ����|       �       �       �           3�     �       �     ��    ���                                                 3�     �       �     ��    `                                                   3�     �            ��    ���                                                 3� (   �       �     ��    (�K                                                3�     �      �     ��                                                       c� 8   �   �   �     ��                                                       8   �   �   �   8   �   �   �   	[refname]       �    :  �         t   @   c� 8   |   �   �    	 ��        	                                               8   |   �   �   8   |   �   �   	[devname]        ����������������    �����       |  ~�{�  ���  }
 �  Switch_Open     Miscellaneous      �?   9 
 ��    h� @T� ��H�}M?0.9m      ��������h�  ��{�G�z�?10m     ��������h� ����      �?0.5     ��������h� ����    ��.A1meg     �������� 45 :�     4       ����4����                        ��xX2_switch_timeX2_switch_time
 9 V            �xSwitches   Generic   X2X2          ��������time controlled switch   TIME_SWITCH�.subckt tswitch 4 5
S 4  5  3 0 switch
V0 3  0 DC 0 PWL ( 0 0
+ {time_on-.000000001} 0
+ {time_on+.000000001}  1
+ {time_off-.000000001} 1
+ {time_off+.000000001} 0)

IVm0 3  0 0

.model switch SW  vt = .5   vh = 0   ron = {res_on}   roff = {res_off}  
.ends   ��     time the switch closes   ParamSubtime_ons              ��    1time the switch opens   ParamSubtime_offs             ��    1resistance when switch closed   ParamSubres_onOhm             ��    1megresistance when switch open   ParamSubres_offOhm               X <�    ����SW+4      PASASW+������<�   ����SW-5      PASASW-   �����SwitchesTime Controlled SwitchGeneric              12 �      �       �   �  �      �   �  �              	voltmeter�        �3 ��    ~           M+i  �   �   �     M-j   �  �          IV_VL    
 1�                   ��                                                           `   M+1�                   ��                                                      �   `   M-3�     `       `     ��    ��                                                3� �   `   �   `     ��                                                        3�    L      \     ��    ��                                                3�     T      T     ��    p�H                                                3� �   X   �   X     ��               	FIXED_ROT                                        a�     <   �   �                   ����                                             <   �   �   c� (   D   �   x     ��                                                      (   D   �   x   (   D   �   x   [value]       X  l  �	  �  (   D   �   x   c�        �   0    	 ��        	                                                      �   0          �   0   	[refname]       @  �  ^	  o         �   0    �  �����  ���      �
     	voltmeter    voltmeter_smallMiscellaneous      �?       f�     h� ����    ���?325.37m      �������� M+M- :�     M+        ����M+����                        ��:�    M-      ����M-����                        ��	voltmeter	voltmeter   _            ��Analog Meters   Generic   IV_VLIV_VL          ����  IVm <�    ����M+M+      PASAM+    ����<�   ����M-M-      PASAM-    ����Analog Meters Generic              12 �  :�    C-      ����C-����                        ���:�    M-      ����M-����                        ��� � 12   12 �     �.    
  �	   "�9    �   �	  �	   � 	      �     	              �   M+0  �   �   �  �   M-1    
   	          VA_IL    	 1�                   ��                                                           @   M+1�                   ��                                                      �   @   M-3� �   @   �   @     ��    ��                                                3�     @       @     ��                                                        3� 4   X   `   X     ��    ��                                                a�        �   d                   ����                                                �   d   �� ����������������  ��          @ @                                           ��d   X    IX1.��X   P        ��X   `    0000@ @ c� $   $   �   L     ��                                                      $   $   �   L   $   $   �   L   [value]       �
  l	  q  �	  $   $   �   L   c�     �����        ��                                                           �����          �����      	[refname]       �
  �  �  �	      �����       �  ���  �  ���  �	     Ammeter    Ammeter_smallMiscellaneous      �?       ��     h� '�     �N$�> 5.99u      �������� M+M- :�     M+        ����M+����                        ���AmmeterAmmeter   �            ��Analog Meters   Generic   VA_ILVA_IL          ����  VAm <�    ����M+M+      PASAM+0�M����<�   ����M-M-      PASAM- ������Analog MetersAmmeterGeneric              11  :�    L-      ����L-����                        ���	 11 	  11 �     �   �  �	   "�;    �   �  �	   �        �                   �   L+K  �   �  �  �   L-L   �   	          L1     1�                    ��                                                           @   L+1�                   ��                                                      �   @   L-�� h   ,   �   T    
                                                           h   ,   �   T   h   ,   �   T   �   @   h   @           �� P   ,   h   T    	                                                           P   ,   h   T   P   ,   h   T   h   @   P   @           �� 8   ,   P   T                                                               8   ,   P   T   8   ,   P   T   P   @   8   @           ��     ,   8   T                                                                   ,   8   T       ,   8   T   8   @       @           3� $   P      X     ��    ��                                                3�    H   $   P     ��     �                                                  3�     P   $   P     ��    ��                                                3�     @       @     ��    p�H	                                                3� �   @   �   @     ��       
                                                c�     \   �   |     ��                                                           \   �   |       \   �   |   [Inductance]       �  
  �  �
      \   �   |   c�         �   $     ��                                                               �   $           �   $   	[refname]       �   	  R  �	          �   $    ���  �  �  �  ���  �  �  �  �     Inductor     Miscellaneous      �?    
   ��  CInductorBehavior     h� ��� �������?100m      ��������h� ���� x     �������� L+L- :�     L+        ����L+����                        ��� Inductor  
              ��Passive   Generic   L1L1          ����  L <�    ����L+L+      PASAL+������<�   ����L-L-      PASAL-P������PassiveInductorGeneric              5  :�     R+        ����R+����                        ��� 5    5  �    �   �  �   R+  �   �       �   R-       	         R     1�                    ��                                                       �   @   R+1�                   ��                                                          @   R-3�    @   $   0     ��    ��)                                                3� 0   P   $   0     ��                                                        3� 0   P   <   0     ��    ��)                                                3� H   P   <   0     ��    p�Z                                                3� H   P   T   0     ��                                                       3� `   P   h   @     ��    D�Z                                                3� �   @   h   @     ��    ��d                                                3� `   P   T   0    	 ��    |�f	                                                3�    @       @    
 ��    <�b
                                                c�     `   �   �     ��                                                           `   �   �       `   �   �   [resistance]           
  �  �
      `   �   �   c�         t   $     ��                                                               t   $           t   $   	[refname]           	  P  �	          t   $    �������������   resistor    resistor DINMiscellaneous      �?       ��  CResistorBehavior     h� �������(\��?0.58      ��������h� ���� 27     ��������h� ����       ��������h� ����       �������� R+R- �:�    R-      ����R-����                        �� resistor                ��Passive   Generic   RR          ����    R <�    ����R+R+      PASAR+JV1.����<�   ����R-R-      PASAR-�)����Passivedefault resistor, 1KGeneric              3 3�t  :�     C+        ����C+����                        ����� J 3   3  �    �   �  �   C-�  �   �        �   C+�   @  �          C1     1�                   ��                                                       �   @   C-1�                   ��                                                          @   C+3�     @   @   @      ��    ���                                                 3� @       @   `     ��    �b�                                                3� `       `   `     ��    ���                                                 3� `   @   �   @     ��    (�K                                                c�     `   �   �     ��                                                           `   �   �       `   �   �   [capacitance]       @  �  �  .	      `   �   �   c�         �   $     ��                                                               �   $           �   $   	[refname]       @  �  �  +          �   $    �����    �      ��     	Capacitor     Miscellaneous      �?       ��  CCapacitorBehavior     h� '  �dy���=20p      ��������h� ���� x     ��������h� ����       ��������h� ����       �������� C+C- �� 	capacitor                ��Passive   Generic   C1C1          ����  C <�    ����C+C+      PASAC+�R����<�   ����C-C-      PASAC-P�����Passive Generic              ?   �C                           . s   G � 2o �        A 
 E 0 q  � = # =                                                     / - w � � W + � � S  � e6{ � U % ' O � ) � � K � Q M � } �� �# R . R   $                           � �  ��      ~ (   �   P         v   �     J     !   � �        0 7d. x � � T � fX z �   N   � * � � � L V & , 5R � � | �    ��  CLetter    �Los dos interruptores se ponen en ON al mismo tiempo.
X2 se pone en OFF, deja de fluir corriente desde la fuente.
X3 sigue en ON, por donde circula la corriente adem�s de por D2.
X3 passa a OFF, entonces la corriente retorna a la fuente a trav�s de D1 y D2.
�   2  �  S  -����Arial����                       Arial            
 h�@ ����        ��������h�             0     ��������h� ����      @5     ��������h�  ʚ;�������?.1     ��������h�@ ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ���� true
     ��������h� ����  false     ��������               
                  h� ����        ��������h� ����       ��������h�  ����       ��������h�@ ����       ��������h�@ ����       ��������               
                  h� ����        ��������h� ����       ��������h�@ ����       ��������h�  ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������               
                 h� ����dec     ��������h� ����     @�@1k     ��������h� ����    ��.A1meg     ��������h� ����       20     ��������h� ���� true     ��������h� ���� true     ��������h� ���� true	     ��������h� ����  false
     ��������               
                 h�  ����        ��������h�  ����       ��������h�  ����       ��������h� ����dec     ��������h� ����       ��������h� ����       ��������h� ����  	     ��������h� ����  
     ��������               
                  	 h� ����        ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������               
                 h� ����        ��������h� ����       ��������h� ����       ��������h� ����dec     ��������h� ����       ��������               
                    h�             0      ��������h�  ��{�G�z�?20m     ��������h� �� �h㈵��>0.01m     ��������h� �� �h㈵��>0.01m     ��������h� ���� True     ��������h� ����  F     ��������h� ���� true     ��������h� ����  false     ��������               
                 h� ����     @�@1K      ��������h�  ����       ��������h�  ����       ��������h�  ����       ��������               
         ��              h�  ����        ��������              
                  h�  ����        ��������              
                                  
                 h�@ ����        ��������h�@ ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ���� true	     ��������h� ����  false
     ��������h� ���� true     ��������h� ����  false     ��������               
                 h� ����       5      ��������h� ����       5     ��������h� ����       5     ��������h� ����       5     ��������h� ����       ��������h� ����  	     ��������h� ����  
     ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ���� true     ��������h�@ ����       ��������h�@ ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����dec     ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ���� true     ��������h� ���� true     ��������h� ���� true     ��������h� ����  false     ��������h� ���� true     ��������h� ����  false      ��������h� ���� true!     ��������h� ����  false"     ��������               
                        h� ����       5      ��������h� ����       5     ��������h� ����       5     ��������h� ����       5     ��������h� ����       ��������h� ����  	     ��������h� ����  
     ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ���� true     ��������h�@ ����       ��������h�@ ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����dec     ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ���� true     ��������h� ���� true     ��������h� ���� true     ��������h� ����  false     ��������h� ���� true     ��������h� ����  false      ��������h� ���� true!     ��������h� ����  false"     ��������               
                 h� ����       5      ��������h� ����       5     ��������h� ����       5     ��������h� ����       5     ��������h� ����       ��������h� ����  	     ��������h� ����  
     ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ���� true     ��������h�@ ����       ��������h�@ ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����dec     ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ���� true     ��������h� ���� true     ��������h� ���� true     ��������h� ����  false     ��������h� ���� true     ��������h� ����  false      ��������h� ���� true!     ��������h� ����  false"     ��������               
                 h� ����       5      ��������h� ����       5     ��������h� ����       5     ��������h� ����       5     ��������h� ����       ��������h� ����  	     ��������h� ����  
     ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ���� true     ��������h�@ ����       ��������h�@ ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����dec     ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ���� true     ��������h� ���� true     ��������h� ���� true     ��������h� ����  false     ��������h� ���� true     ��������h� ����  false      ��������h� ���� true!     ��������h� ����  false"     ��������               
                 h�@ ����        ��������h�@ ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����decade     ��������h� ���� true     ��������h� ���� true     ��������h� ���� true     ��������h� ����  false     ��������               
                 h� ����        ��������h� ����       ��������h�@ ����       ��������h�  ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������h� ����       ��������               
                        h� ����dec     ��������h� ����     @�@1k     ��������h� ����    ��.A1meg     ��������h� ����       20     ��������h� ����        0     ��������h� ����        0     ��������h� ���� true	     ��������h� ���� true
     ��������h� ����      I@50     ��������h� ���� true     ��������h� ����  false     ��������               
                         / h� ���� x'     ��������h�     �-���q=1E-12     ��������h� @B -C��6?1E-4     ��������h� ���� x     ��������h� ���� x     ��������h� ���� x     ��������h� ���� x     ��������h� ���� x     ��������h� ���� x     ��������h� ���� x	     ��������h� ���� x!     ��������h� ����    �  500
     ��������h� ���� x     ��������h� ����    �  500     ��������h� ���� x$     ��������h� ���� x$     ��������h� ���� x%     ��������h� ���� x"     ��������h�  ���� x*     ��������h� ���� x     ��������h� ���� x     ��������h� ���� x     ��������h� ���� x&     ��������h� ���� x     ��������h� ���� x     ��������h� ���� x     ��������h� ���� x+     ��������h� ���� x,     ��������h� ���� x-     ��������h� ���� xg     ��������h� ���� xf     ��������h� ���� xd     ��������h� ���� xe     ��������h� ���� xh     ��������h� ���� xj     ��������h� ���� xi     ��������h� ���� xk     ��������h� ����    e��A1Gl     ��������h�             0�     ��������h� ����      @5�     ��������h� ����      @2.5�     ��������h� ����      �?.5�     ��������h� ����      @4.5�     ��������h� 
   ��&�.>1n�     ��������h� 
   ��&�.>1n�     ��������h� 
   ��&�.>1n�     ��������h� 
   ��&�.>1n�     ��������           ��  CPrimitiveModel    d1n4007   h�    1�a��%>2.55e-9      ��������h� ���� 27     ��������h�  �/�$��?0.042     ��������h� ����      �?1.75     ��������h�  �  ��v��(�>5.76e-6     ��������h�     �]}IW�=1.85e-11     ��������h� ����      �?0.75     ��������h� ����Zd;�O�?0.333     ��������h� ���� 1.11	     ��������h� ���� 3.0
     ��������h�      0     ��������h� ���� 1     ��������h� ���� 0.5     ��������h� ����     @�@1000     ��������h� � Ǯ���?9.86e-5     ��������     Diode Generic��   CPrimitiveModelType Junction Diode model����DD   ������ 1.0E-14Saturation current    ProcessisAmp0       e     ������ 27!Parameter measurement temperature    ProcesstnomDeg C0     s     ������ 0Ohmic resistance    ProcessrsOhm0      f     ������ 1Emission Coefficient    Processn 0      g     ������ 0Transit Time    Processttsec0     h     ������ 0Junction capacitance    ProcesscjoF0     i     ������ 0     Processcj0F0     i     ������ 1Junction potential    ProcessvjV0      j     ������ 0.5Grading coefficient    Processm 0      k     ������ 1.11Activation energy    ProcessegeV0     	 l     ������ 3.0#Saturation current temperature exp.    Processxti 0     
 m     ������ 0flicker noise coefficient    Processkf 0      t     ������ 1flicker noise exponent    Processaf 0      u     ������ 0.5#Forward bias junction fit parameter    Processfc 0      n     ������ infReverse breakdown voltage    ProcessbvV0      o     ������ 1.0e-3$Current at reverse breakdown voltage    ProcessibvA0      p     ������  Ohmic conductance    ProcesscondMho     r        D��     &� �                Ariald     h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  COpAnal                         
                        ����            
G3                ��  TSignal                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                      v(iv_vl)       ����                  B�                     	i(va_ix1)       ����                  B�                     i(va_il)       ����                  B�                      	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CDCsweep       
 	
               
                       ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                       v(iv_vl)       ����                  B�                      	i(va_ix1)       ����                  B�                      i(va_il)       ����                  B�                       	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACsweep        !"#$%&'(               
                       ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                      v(iv_vl)       ����                  B�                     	i(va_ix1)       ����                  B�                     i(va_il)       ����                  B�                      	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  �� 
 CTranSweep       ?@ABCDEF               
                       ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                       v(iv_vl)       ����                  B�                      	i(va_ix1)       ����                  B�                      i(va_il)       ����                  B�                       	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACdisto        :;<=>               
                           ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                       v(iv_vl)       ����                  B�                      	i(va_ix1)       ����                  B�                      i(va_il)       ����                  B�                       	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��        h� ����        ��������h� ����       ��������h� ����       ��������h� ����dec     ��������h� ����       ��������               
                          ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                       v(iv_vl)       ����                  B�                      	i(va_ix1)       ����                  B�                      i(va_il)       ����                  B�                       	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��        h� ����        ��������h� ����       ��������h� ����       ��������h� ����dec     ��������h� ����       ��������               
                          ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                       v(iv_vl)       ����                  B�                      	i(va_ix1)       ����                  B�                      i(va_il)       ����                  B�                       	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��        h� ����        ��������h� ����       ��������h� ����       ��������h� ����dec     ��������h� ����       ��������               
                           ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                       v(iv_vl)       ����                  B�                      	i(va_ix1)       ����                  B�                      i(va_il)       ����                  B�                       	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��        h� ����        ��������h� ����       ��������h� ����       ��������h� ����dec     ��������h� ����       ��������               
                          ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                       v(iv_vl)       ����                  B�                      	i(va_ix1)       ����                  B�                      i(va_il)       ����                  B�                       	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��        h� ����        ��������h� ����       ��������h� ����       ��������h� ����dec     ��������h� ����       ��������               
         �             	    ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                       v(iv_vl)       ����                  B�                      	i(va_ix1)       ����                  B�                      i(va_il)       ����                  B�                       	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACnoise        )*+,-./0               
                    
    ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                      v(iv_vl)       ����                  B�                     	i(va_ix1)       ����                  B�                     i(va_il)       ����                  B�                      	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��         h�  ����        ��������h�  ����       ��������h�  ����       ��������h� ����dec     ��������h� ����       ��������h� ����       ��������h� ����  	     ��������h� ����  
     ��������              
                        ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                      v(iv_vl)       ����                  B�                     	i(va_ix1)       ����                  B�                     i(va_il)       ����                  B�                      	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CFourier        GHIJ               
         ��                   ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                      v(iv_vl)       ����                  B�                     	i(va_ix1)       ����                  B�                     i(va_il)       ����                  B�                      	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACpz        	 123456789               
                       ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                      v(iv_vl)       ����                  B�                     	i(va_ix1)       ����                  B�                     i(va_il)       ����                  B�                      	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CDCtf                        
                       ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                      v(iv_vl)       ����                  B�                     	i(va_ix1)       ����                  B�                     i(va_il)       ����                  B�                      	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CDCsens                         
                       ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                       v(iv_vl)       ����                  B�                      	i(va_ix1)       ����                  B�                      i(va_il)       ����                  B�                       	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j                  ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                      v(iv_vl)       ����                  B�                     	i(va_ix1)       ����                  B�                     i(va_il)       ����                  B�                      	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CShow         K              
                       ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                      v(iv_vl)       ����                  B�                     	i(va_ix1)       ����                  B�                     i(va_il)       ����                  B�                      	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CShowmod         L              
                       ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                      v(iv_vl)       ����                  B�                     	i(va_ix1)       ����                  B�                     i(va_il)       ����                  B�                      	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  �� 
 CLinearize        h�  ����        ��������               
                       ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                      v(iv_vl)       ����                  B�                     	i(va_ix1)       ����                  B�                     i(va_il)       ����                  B�                      	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CParamTranSweep        MNOPQRSTUVWXY               
                       ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                      v(iv_vl)       ����                  B�                     	i(va_ix1)       ����                  B�                     i(va_il)       ����                  B�                      	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  S              ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                       v(iv_vl)       ����                  B�                      	i(va_ix1)       ����                  B�                      i(va_il)       ����                  B�                       	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CParamACSweep        �������������               
                       ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                      v(iv_vl)       ����                  B�                     	i(va_ix1)       ����                  B�                     i(va_il)       ����                  B�                      	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CMonteCarlo_op        Z[\]^_`abcdefghijklmnopqrstu               
                              ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                      v(iv_vl)       ����                  B�                     	i(va_ix1)       ����                  B�                     i(va_il)       ����                  B�                      	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CMonteCarlo_dc        vwxyz{|}~������������������               
                       ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                       v(iv_vl)       ����                  B�                      	i(va_ix1)       ����                  B�                      i(va_il)       ����                  B�                       	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CMonteCarlo_ac        ����������������������������               
                       ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                      v(iv_vl)       ����                  B�                     	i(va_ix1)       ����                  B�                     i(va_il)       ����                  B�                      	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CMonteCarlo_tran        ����������������������������               
                       ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                       v(iv_vl)       ����                  B�                      	i(va_ix1)       ����                  B�                      i(va_il)       ����                  B�                       	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACsens        �����������               
                              ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                       v(iv_vl)       ����                  B�                      	i(va_ix1)       ����                  B�                      i(va_il)       ����                  B�                       	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CNetworkAnalysis        �����������               
                       ����            P               B�                        v(13)       ����                  B�                       v(3)       ����                  B�                       v(4)       ����                  B�                       v(5)       ����                  B�                       v(9)       ����                  B�                       v(7)       ����                  B�                       v(8)       ����                  B�                       v(10)       ����                  B�                       v(11)       ����                  B�	                       v(12)       ����                  B�
                       v(iv_vl)       ����                  B�                      	i(va_ix1)       ����                  B�                      i(va_il)       ����                  B�                       	v(iv_vx1)       ����                  B�                       i(x2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j                  ����            P              33�=           ��   CDigSimResTemplate                ���       ����  ����:�0�yU>20.00n���   ����                       Arial����                       Arial����                       Arial  �   �  �                                ����  ���� ������       ����  ���� ������                 �               ����  �����       200������         0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial      �       �         �     �   �  �  Circuit1                  ����  ��    ��������                                                                                                                                                                         g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     ��   CPackageAliasSuperPCBStandardDIODE3      H�Eagle	DIODE.LBRDO41-7   AC  H�Orcad 	DAX2/DO41      H�	Ultiboard	L7DIO.l55DIO_DO41              A      g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     H�SuperPCBStandardDIODE3      H�Eagle	DIODE.LBRDO41-7   AC  H�Orcad 	DAX2/DO41      H�	Ultiboard	L7DIO.l55DIO_DO41              A                                              �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                      �  �                a�         �  @                  ���                                                  �  @  3�     <   �  <     ��                                                        3�     |   �  |     ��                                                        3�     �   �  �     ��                                                        3�     �   �  �     ��                                                        c� �      �  4     ��                                                      �      �  4   �      �  4   [title]                                       c� �   D   �  t     ��                                                      �   D   �  t   �   D   �  t   [description]                                       c� `   �   h  �     ��                                                      `   �   h  �   `   �   h  �   [id]                                       c� �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       c�      �   8    ��        	                                                   �   8       �   8  Date :       �    8
  �                  c� �     �  4   	 ��        
                                              �     �  4  �     �  4  [date]                                       c�       t   8    
 ��                                                            t   8         t   8   Title :       �    
  �                  c�    L   �   x     ��                                                         L   �   x      L   �   x   Description :       �  �  �  �                  c�    �   �   �     ��                                                         �   �   �      �   �   �   ID :       �  �  �	  T                  c�    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �  L  (                     STUVWXYZ[]^_`a          \     	title box    Analog Misc      �?    9 
 ��     h�  ����        ��������h�  ����       ��������h�  ����       ��������h�  ����       ��������h�  ����       ��������        9                                      �������� ����     ��            title                ��            description               ��            id               ��            designer               ��            date                           ����            `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                                                                                            2         �  �              � � �                   ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                          �   ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    
cgs 76         47 80moh5.6 (�P    mvrd nmodel ��P�P      B�                      TIME� # ) time                      B�                        v(3)      v(3)    TIME                 B�                      	i(va_ix1)�   � 	i(va_ix1)    TIME                 B�    (v(7)-v(3))                   v(IV_VL)� �   v(IV_VL)    TIME                 B�                      i(va_il)  � � i(va_il)    TIME                 B�    v(5)                   	v(IV_Vx1)� �   	v(IV_Vx1)    TIME                 B�    v(iv_vx1)*i(va_ix1)                    Pin� # )  ����TIME                 B�                        v(5)      v(5)    TIME                 B�                      i(va_d2)    � i(va_d2)    TIME                 B�                      i(va_x2)� �   i(va_x2)    TIME                 B�                      i(va_x1)�   � i(va_x1)    TIME                 B�                      i(va_d1)  � @ i(va_d1)    TIME                 B�                        v(7)      v(7)    TIME                           2         �  �           Time  � � �              �     ����                       Arial����                       Arial                              ����  ����ё�[W?1.425662e-003����       ����  ����� �6lD?6.109980e-004��;]       ����  �������հ	@3.211344e+000������      ����  ������>��Nڿ-4.110512e-001������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 1m  0                            100   100                                                             1m  0                            100   100                                1m  0                            100   100                                1m  0                            100   100                                                 
                 1m  0                            100   100                            ��   CPartPackage     ��   CPackageg   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     MNOP   }��/� �g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     IJKL      ��   CMiniPartPin    ����C+C+     PASC+�      ��   ����C-C-     PASC-�     capacitor_genericcapacitor_generic                          ��    ����11     PAS1�      ��   ����22     PAS2�     BatteryBattery                          ��    ����R+R+     PASR+      ��   ����R-R-     PASR-     RR                          ��    ����GndGnd     GNDGnd}      GndGnd                  ��    ����M+M+     PASM+i      ��   ����M-M-     PASM-j     	voltmeter	voltmeter                          ��    ����M+M+     PASM+2      ��   ����M-M-     PASM-3     Ammeter2Ammeter2                          ��    ����M+M+     PASM+2      ��   ����M-M-     PASM-3     Ammeter2Ammeter2                          ��    ����M+M+     PASM+2      ��   ����M-M-     PASM-3     Ammeter2Ammeter2                          ��    ����SW+4     PASSW+=      ��   ����SW-5     PASSW->     switch_timeswitch_time                          ��    ����L+L+     PASL+K      ��   ����L-L-     PASL-L     InductorInductor                          ��    ����M+M+     PASM+0      ��   ����M-M-     PASM-1     AmmeterAmmeter                          ��    ����M+M+     PASM+k      ��   ����M-M-     PASM-l     
Voltmeter2
Voltmeter2                       � ��    ����D+D+     PASA       ��   ����D-D-     PASK       �   ��   CPackagePin 1 D+PAS  AA�� 2 D-PAS  AKDiodeDiode	Fairchild      1n4007 D1n4007D2            diode-21n40071n4007                       ~ ��    ����D+D+     PASA       ��   ����D-D-     PASK       2  �� 1 D+PAS  AA�� 2 D-PAS  AKDiodeDiode	Fairchild      1n4007 D1n4007D1            diode-21n40071n4007                          ��    ����M+M+     PASM+2      ��   ����M-M-     PASM-3     Ammeter2Ammeter2                          ��    ����M+M+     PASM+2      ��   ����M-M-     PASM-3     Ammeter2Ammeter2                          ��    ����SW+4     PASSW+=      ��   ����SW-5     PASSW->     switch_timeswitch_time                                                                                                                                                                                         ��    �Z�P��,�                        ��                                                                                                            (f    x=f � �'f                           �(f                            ,�e    �f � ��e                           ��e                                     �  � ���� �                         .I                                                                                                        
                                                                                                                             |                               �     � �� �� (�K                        �                              ��    ��������P��                        ��                            �V�    (W�`W��W��W�                        �Y�                            Їl    `�l(�l`-j �W                         �W                            t�@
    L �k��
>ENDDATA
                        
JV1                            p�<        ��<x�                           �                            \       |     ��                                                              �a�    �E��E�@F�xF�                        �o�                                         �rP��                                 2 2 2 2 d                                                                   