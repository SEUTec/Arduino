    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz    ��  CPart    �����   �  �  �����   �  �              voltage_source��  CIntPin    ��  CWire     �        �       �      @      �      @              BUZ11 �   �     �    
     �           �   �           �   �               Gnd ��  CExtPin    ��  CVertex   �  @   ��  CSegment
   �   �  `	                 �   �   �  @   �   �   �  �
                  �   �   �  @   �   �   �  �                                       �    �(   @  @   �   �%   @  `	                  �    �#      @     �   �&      �
   "         !                                   `       Gnd}   `  @          gnd1     ��   CPin                    ��                                                               Gnd��  TLine                   ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        &�         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        &�    ,   4   ,     ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        &�    8   (   8     ��    p�Z         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         % ' ( *   )      Ground    
Ground DINMiscellaneous      �?       ��   CGroundBehavior       Gnd ��   CBehPin     Gnd        ����Gnd����                        ��gndgnd                 . Analog Meters   Generic   gnd1gnd1          ����  gnd ��   CPartPin    ����GndGnd      GNDAGnd �)����SourcesGroundGeneric              0 	 �   
     0 �   
    �           �   �          �   �              Battery�    �    4 �    5    �       _   @  �      _   @  �              Ammeter26 �   �    8 �   9   �       �      @      �      @              BUZ11�    �    < �    =    �   �����   �  �  �����   �  �              voltage_source> �   �    �    A    �       �   �  �       �   �  �               RB �   �    �   E    3 D �   E   �	       �      @      �      @              BUZ11�    �    I �    J    �
   �����   �  �  �����   �  �              voltage_sourceK �   E   L 3 �    �    �      �   �"   �  �   P �   Q �   �  �   R    	             O        
               V+ ����   �!   �  �   �	   U �
   �  �   �   �   �      X    	    W     V �   W �   �  �   Z             �   W �   �      �   ] �   �      ^            \ �   ] �   �  �   `                               
          �  V-��R �            V3     $�                   ��                                                           `   V+$�                   ��                                                          �   V-��  TEllipse     �   �����                   ����                                         �����       �   �����       �   &�    �   �����     ��     �                                                 &�     �       �     ��                                                        &�     �       �     ��                                                        &�     \       �     ��                                                        &� �����   
   �    
 ��                	FIXED_ROT                                        ��  
 TTextField \   `   \   `     ��                                                      \   `   \   `   \   `   \   `           �     �                   k� 0   �   �   �     ��        	                                               0   �   �   �   0   �   �   �   [dc]       p  �  �  F          p   @   k� 0   \   �   �    	 ��        
                                               0   \   �   �   0   \   �   �   	[refname]       p    �  �      ����t       e   f g i c h l m n       j     b  �  Voltage Source    Voltage Source DINRoot      �?       ��  CVSourceBehavior     ��  CValue ����        0      ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       �������� V+V- -�     V+        ����V+����                        ��-�    V-      ����V-����                        ��volt_sourcevolt_source   +0            ~  Sources   Generic   V3V3          ����       q�0����      @5      ��������q�0            0     ��������q�0            0     ��������q�0�� �h㈵��>10u     ��������q�0P�  �h㈵��>5u     ��������q�0���{�G�zt?5m     ��������q�0 ��{�G�z�?10m     ��������    q�0            0      ��������q�0����      @5     ��������q�0����     ��@10k     ��������q�0            0     ��������q�0            0     ��������    q�0            0      ��������q�0����      �?1     ��������q�0����      �?1     ��������q�0            0     ��������q�0����      �?1     ��������    q�0            0      ��������q�0����      �?1     ��������q�0            0     ��������q�0 N  �����>2u     ��������q�0'  ���ư>1u     ��������q�0'  ���ư>1u     ��������    q�  ���� 0 0      ��������                0      �������� ����       �������� ����       �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������               V /�    ����V+V+      PWR+AV+�eW����/�   ����V-V-      PWR-AV-�3W����Sources Generic              9  -�     1       ����gate����                        ��~  9   H 9 G �   9   H 7 �    S        �  Gate@
G�   �   �  �   �   �   �  �   �   �   @  �   �   � �   @  �   �            �     �     �   �   �  �   �        �     �     �        	         �   Drain�r�?�   Y      @  SourceE�@ �  �          X4     $�                    ��                                                           �   Gate$�                   ��                                                      `   @   Drain$�                   ��                                                      `   �   Source&�     �   ,   �     ��                                                        &� ,   d   ,   �     ��                                                        &� 8   T   8   l     ��                                                        &� 8   `   `   `     ��                                                        &� `   @   `   `     ��                                                        &� 8   �   `   �     ��                                                        &� `   �   `   �    	 ��        	                                                &� D   �   P   �    
 ��        
                                                &� P   t   D   �     ��                                                        &� 8   �   `   �     ��                                                        &� `   �   `   �     ��                                                        &� 8   x   8   �     ��                                                        &� 8   �   8   �     ��                                                        k� ����   �   <     ��                                                       ����   �   <   ����   �   <   	[refname]       �  (    �  ����   �   <   k� ���������        ��                                                       ���������      ���������      	[devname]        �������������������������       � � � � � � � � � � � � � � � � �   �      
Mos 3 nmos     Miscellaneous      �?   #    X /�    ����Gate1      PASAGate   �����/�   ����Source2      PASASource rel����/�   ����Drain3      PASADrain�����MOSFETsMOSFETsSiemensTO-220             3 M �    E    �       �   �  �      �   �  �              	voltmeter� �   A   � 6 �    [           M+    �   �   �
  �   �   � �   @  �   �   �    @      �        �     � �   � �      �   �            �   � �	   @      �   �    
      �         �     � �   � �$   @  �   �                                     �     M-    �  �          IVm1    
 $�                   ��                                                           `   M+$�                   ��                                                      �   `   M-&�     `       `     ��    ��                                                &� �   `   �   `     ��                                                        &�    L      \     ��    ��                                                &�     T      T     ��    p�H                                                &� �   X   �   X     ��               	FIXED_ROT                                        �� 
 TRectangle     <   �   �                   ����                                             <   �   �   k� (   D   �   x     ��                                                      (   D   �   x   (   D   �   x   [value]       X  L  0	  �  (   D   �   x   k�        �   0    	 ��        	                                                      �   0          �   0   	[refname]       @  �  0	  D         �   0    �   � � � � �   � � �       � 
     	voltmeter    voltmeter_smallMiscellaneous      �?       ��   CVoltmeterBehavior     q� ����  ���-@ 5.04      �������� M+M- -� 4  M+        �  M+����                        ��-� 4  M-      �  M-����                        ��	voltmeter	voltmeter   _            � � Analog Meters   Generic   IVm1IVm1          ����  IVm /�    ����M+M+      PASAM+� �
    /�   ����M-M-      PASAM-       Analog Meters Generic              3  -�    3      ����drain����                        ��-�    R-      ����R-����                        ��� -�    2      ����source����                        ��  3  C 3 �    �    �  �   R+  �   _       �   R-   �  `         RL     $�                    ��                                                       �   @   R+$�                   ��                                                          @   R-&�    @   $   0     ��    ��)                                                &� 0   P   $   0     ��                                                        &� 0   P   <   0     ��    ��)                                                &� H   P   <   0     ��    p�Z                                                &� H   P   T   0     ��                                                       &� `   P   h   @     ��    D�Z                                                &� �   @   h   @     ��    ��d                                                &� `   P   T   0    	 ��    |�f	                                                &�    @       @    
 ��    <�b
                                                k�     `   �   �     ��                                                           `   �   �       `   �   �   [resistance]       �  �  	        `   �   �   k�         t   $     ��                                                               t   $           t   $   	[refname]       �  `   	             t   $    � � � � � � � � � � � � �    resistor    resistor DINMiscellaneous      �?       ��  CResistorBehavior     q� ����      6@22      ��������q� ���� 27     ��������q� ����       ��������q� ����       �������� R+R- -�     R+        ����R+����                        ���  resistor                � � Passive   Generic   RLRL          ����    R /�    ����R+R+      PASAR+�)����/�   ����R-R-      PASAR-JV1.����Passivedefault resistor, 1KGeneric              6 �   A   ; 6 � @ �   A   �       �      @      �      @              BUZ11�    �    � �        �   �����   �  �  �����   �  �              voltage_source�   
    0 �    �'      `	   �!   �*       	   �   �   `   	                                         V+@
G�   #       �  V-�@
    @         V4     $�                   ��                                                           `   V+$�                   ��                                                          �   V-d�     �   �����                   ����                                         �����       �   �����       �   &�    �   �����     ��                                                        &�     �       �     ��                                                        &�     �       �     ��                                                        &�     \       �     ��    ��V                                                &� �����   
   �    
 ��                	FIXED_ROT                                        k� \   `   \   `     ��                                                      \   `   \   `   \   `   \   `           4  `	  4  `	                k� 0   �   �   �     ��        	                                               0   �   �   �   0   �   �   �   [dc]       �  �	  �  �
          p   @   k� 0   \   �   �    	 ��        
                                               0   \   �   �   0   \   �   �   	[refname]       �  T	  0  �	      ����t                    �  Voltage Source    Voltage Source DINRoot      �?       o�     q� ����        0      ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       �������� V+V- -�     V+        ����V+����                        ��-�    V-      ����V-����                        ��volt_sourcevolt_source   +0            #$Sources   Generic   V4V4          ����       q�0����      @5      ��������q�0            0     ��������q�0            0     ��������q�0�� �h㈵��>10u     ��������q�0P�  �h㈵��>5u     ��������q�0���{�G�zt?5m     ��������q�0 ��{�G�z�?10m     ��������    q�0            0      ��������q�0����      @5     ��������q�0����     ��@10k     ��������q�0            0     ��������q�0            0     ��������    q�0            0      ��������q�0����      �?1     ��������q�0����      �?1     ��������q�0            0     ��������q�0����      �?1     ��������    q�0            0      ��������q�0����      �?1     ��������q�0            0     ��������q�0 N  �����>2u     ��������q�0'  ���ư>1u     ��������q�0'  ���ư>1u     ��������    q�  ���� 0 0      ��������                0      �������� ����       �������� ����       �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������               V /�    ����V+V+      PWR+AV+�B<
����/�   ����V-V-      PWR-AV-DATA����Sources Generic              10  � # 10   � 10 �   
    � 0 � �    	      �  Gate.I ��   �       �   Drain3305�          @  SourceA
>D @            X5     $�                    ��                                                       `   �   Gate$�                   ��                                                          @   Drain$�                   ��                                                          �   Source&� `   �   4   �     ��    ATA
                                                &� 4   d   4   �     ��    5227                                                &� (   T   (   l     ��     �)�                                                &� (   `       `     ��    4�5
                                                &�     @       `     ��     �                                                &� (   �       �     ��    ��@                                                &�     �       �    	 ��    �@
	                                                &�    �      �    
 ��    ATA

                                                &�    t      �     ��    5322                                                &� (   �       �     ��     �
                                                &�     �       �     ��    ���
                                                &� (   x   (   �     ��     ��                                                &� (   �   (   �     ��    ��@                                                k� ����   �   <     ��                                                       ����   �   <   ����   �   <   	[refname]       4  h  �    ����   �   <   k� ���������        ��                                                       ���������      ���������      	[devname]        �������������������������       CDEFGHIJKLMNOPQRT  S     
Mos 3 nmos     Miscellaneous      �?   #    X /�    ����Gate1      PASAGateG7  ����/�   ����Source2      PASASource>
 A����/�   ����Drain3      PASADrainTAB ����MOSFETsMOSFETsSiemensTO-220             6  � � � -�    V-      ����V-����                        ���  6  ? 6 �    �          �    �      �   [�   �   `  �   ]        \        Z                      V+    �   �       �  V-�V              V2     $�                   ��                                                           `   V+$�                   ��                                                          �   V-d�     �   �����                   ����                                         �����       �   �����       �   &�    �   �����     ��     �                                                 &�     �       �     ��     �                                                 &�     �       �     ��     �                                                 &�     \       �     ��     �                                                 &� �����   
   �    
 ��     �         	FIXED_ROT                                        k� \   `   \   `     ��                                                      \   `   \   `   \   `   \   `           4     4                   k� 0   �   �   �     ��        	                                               0   �   �   �   0   �   �   �   [dc]       �  �  �  F          p   @   k� 0   \   �   �    	 ��        
                                               0   \   �   �   0   \   �   �   	[refname]       �    0  �      ����t       b  cdfaehij      g    ` �  Voltage Source    Voltage Source DINRoot      �?       o�     q� ����        0      ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       �������� V+V- -�     V+        ����V+����                        ��Xvolt_sourcevolt_source   +0            xXSources   Generic   V2V2          ����       q�0            0      ��������q�0����      @5     ��������q�0            0     ��������q�0�� �h㈵��>10u     ��������q�0P�  �h㈵��>5u     ��������q�0���{�G�zt?5m     ��������q�0 ��{�G�z�?10m     ��������    q�0            0      ��������q�0����      @5     ��������q�0����     ��@10k     ��������q�0            0     ��������q�0            0     ��������    q�0            0      ��������q�0����      �?1     ��������q�0����      �?1     ��������q�0            0     ��������q�0����      �?1     ��������    q�0            0      ��������q�0����      �?1     ��������q�0            0     ��������q�0 N  �����>2u     ��������q�0'  ���ư>1u     ��������q�0'  ���ư>1u     ��������    q�  ���� 0 0      ��������                0      �������� ����       �������� ����       �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������               V /�    ����V+V+      PWR+AV+5   ����/�   ����V-V-      PWR-AV-03
J����Sources Generic              8  � x 8   ; 8 � : �    ^      �  Gate  �?�   �       �   Drain8�T�   �       @  Source     @  �         X3     $�                    ��                                                       `   �   Gate$�                   ��                                                          @   Drain$�                   ��                                                          �   Source&� `   �   4   �     ��                                                        &� 4   d   4   �     ��                                                        &� (   T   (   l     ��                                                        &� (   `       `     ��                                                        &�     @       `     ��                                                        &� (   �       �     ��                                                        &�     �       �    	 ��        	                                                &�    �      �    
 ��        
                                                &�    t      �     ��                                                        &� (   �       �     ��                                                        &�     �       �     ��                                                        &� (   x   (   �     ��                                                        &� (   �   (   �     ��                                                        k� ����   �   <     ��                                                       ����   �   <   ����   �   <   	[refname]       4  (  �  �  ����   �   <   k� ���������        ��                                                       ���������      ���������      	[devname]        �������������������������       �����������������  �     
Mos 3 nmos     Miscellaneous      �?   #    X /�    ����Gate1      PASAGate   �����/�   ����Source2      PASASource�W����/�   ����Drain3      PASADrain ?X����MOSFETsMOSFETsSiemensTO-220             7 �  -�    M-      ����M-����                        ���  7  7 7 �    �   �      �   ��   �  `   �                       `   �  M+2  �   �   `   `   M-3   @            VA_Ix1    	 $�                    ��                                                           �   M+$�                   ��                                                              M-&�     �       �     ��                                                        &�     <             ��                                                        ր @   <   �����                  ����                                         ����<   @   �   &� ����x   ����L     ��                                                        ��  TPolygon  ������� �������  ��          @ @                                           ��  TPoint����H    ��b������T    
>DA������T    uT@ @ k� ����D   <   |     ��                                                      ����D   <   |   ����D   <   |   [value]         �  �  �     D   �   |   k�    �����        ��                                                          �����         �����      	[refname]       L    �  �     �����      
 ������  ���	   Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       ��   CAmmeterBehavior     q� ����   `���?226.19m      �������� M+M- -�     M+        ����M+����                        ���AmmeterAmmeter   V            ��Analog Meters   Generic   VA_Ix1VA_Ix1          ����  VAm /�    ����M+M+      PASAM+8�W����/�   ����M-M-      PASAM-��W����Analog MetersAmmeter-verticalGeneric              5  -�     1       ����1����                        ��� 5   3 5 2 �    �   `       1�  �      `   �  2�   @  `          X1     $�                    ��                                                               1$�                   ��                                                          �   2&�             $     ��    ��)                                                &�     \       �     ��                                                        &�    8   0   8    	 ��    ��)                                                &�     H   @   H     ��    p�Z                                                &�     $   @   $     ��                                                       &�    \   0   \     ��    D�Z                                                &�               ���                                                      &�               ���   �Z	                                                k� `          $    
 ��        
                                               `          $   `          $   	[devname]        ����������������`          $   k� `   $      H     ��                                                       `   $      H   `   $      H   	[refname]       `  �  �  l  `   $      H    ��������    ��    �  �     Battery     Miscellaneous      �?    9 
 ��  CParamSubBehavior     q� ����      @5      �������� 12 �-�    2      ����2����                        ��BatteryBattery  9 i             ��Sources   Generic   X1X1          ������   CParamSubModelType��    BATTERY2.SUBCKT Xbattery 1 2
V1 1 2 DC {voltage}
.ENDS
   ��  	 CParmDefn    1battery voltage   ParamSubvoltageV                X /�    ����11      PASA10Ab����/�   ����22      PASA2�1b����SourcesBatteryGeneric              0 ? -�    V-      ����V-����                        ��� �. $  0    0 F �    �   �   	   �   �   �   	   �    ��)   �  `	   �             �    �                   �  Gatey  �   a      �   Drainw  �         @  Sourcex   �             X2     $�                    ��                                                           �   Gate$�                   ��                                                      `   @   Drain$�                   ��                                                      `   �   Source&�     �   ,   �     ��    ��)                                                &� ,   d   ,   �     ��                                                       &� 8   T   8   l     ��    ��)                                                &� 8   `   `   `     ��    p�Z                                                &� `   @   `   `     ��                                                       &� 8   �   `   �     ��    �Z                                                &� `   �   `   �    	 ��       	                                                &� D   �   P   �    
 ��        
                                                &� P   t   D   �     ��                                                        &� 8   �   `   �     ��                                                        &� `   �   `   �     ��                                                        &� 8   x   8   �     ��                                                        &� 8   �   8   �     ��                                                        k� ����   �   <     ��                                                       ����   �   <   ����   �   <   	[refname]       �  h      ����   �   <   k� ���������        ��                                                       ���������      ���������      	[devname]        �������������������������       �����������������  �     
Mos 3 nmos     Miscellaneous      �?   #    X /�    ����Gate1      PASAGate    ����/�   ����Source2      PASASource � ����/�   ����Drain3      PASADrain7   ����MOSFETsMOSFETsSiemensTO-220             4  -�     V+        ����V+����                        ���  4    4 1 �    �          V+g  �          �  V-h   �  @         V1     $�                   ��                                                           `   V+$�                   ��                                                          �   V-d�     �   �����                   ����                                         �����       �   �����       �   &�    �   �����     ��    ��)                                                &�     �       �     ��    ��`                                                &�     �       �     ��    ��)                                                &�     \       �     ��    p�Z                                                &� �����   
   �    
 ��               	FIXED_ROT                                        k� \   `   \   `     ��                                                      \   `   \   `   \   `   \   `           �  `	  �  `	                k� 0   �   �   �     ��        	                                               0   �   �   �   0   �   �   �   [dc]         �	  H  �
          p   @   k� 0   \   �   �    	 ��        
                                               0   \   �   �   0   \   �   �   	[refname]         T	  �  �	      ����t          	          � �  Voltage Source    Voltage Source DINRoot      �?       o�     q� ����        0      ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       �������� V+V- ��volt_sourcevolt_source   +0            ��Sources   Generic   V1V1          ����       q�0            0      ��������q�0����      @5     ��������q�0            0     ��������q�0�� �h㈵��>10u     ��������q�0P�  �h㈵��>5u     ��������q�0���{�G�zt?5m     ��������q�0 ��{�G�z�?10m     ��������    q�0            0      ��������q�0����      @5     ��������q�0����     ��@10k     ��������q�0            0     ��������q�0            0     ��������    q�0            0      ��������q�0����      �?1     ��������q�0����      �?1     ��������q�0            0     ��������q�0����      �?1     ��������    q�0            0      ��������q�0����      �?1     ��������q�0            0     ��������q�0 N  �����>2u     ��������q�0'  ���ư>1u     ��������q�0'  ���ư>1u     ��������    q�  ���� 0 0      ��������                0      �������� ����       �������� ����       �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������               V /�    ����V+V+      PWR+AV+NDDA����/�   ����V-V-      PWR-AV- � ����Sources Generic               3 C  � 7 ; ? H L � 	 	 	 
  E 5 A 9 = J  " " " [� "  ^  � � V  ` X �  � � �]� � � \ P R Z   �  �  �+ + + � �   a �	�  � W  ] � _ � � �� [ � � ^� Z\Y � S � O U Q ! �  #  �             
 q�@ ����        ��������q�             0     ��������q� ����      @5     ��������q�  ʚ;�������?.1     ��������q�@ ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ���� true
     ��������q� ����  false     ��������               
                  q� ����        ��������q� ����       ��������q�  ����       ��������q�@ ����       ��������q�@ ����       ��������               
                  q� ����        ��������q� ����       ��������q�@ ����       ��������q�  ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������               
                 q� ����dec     ��������q� ����     @�@1k     ��������q� ����    ��.A1meg     ��������q� ����       20     ��������q� ���� true     ��������q� ���� true     ��������q� ���� true	     ��������q� ����  false
     ��������               
                 q�  ����        ��������q�  ����       ��������q�  ����       ��������q� ����dec     ��������q� ����       ��������q� ����       ��������q� ����  	     ��������q� ����  
     ��������               
                  	 q� ����        ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������               
                 q� ����        ��������q� ����       ��������q� ����       ��������q� ����dec     ��������q� ����       ��������               
                    q�             0      ��������q�  ��{�G�z�?20m     ��������q� @B -C��6?0.1m     ��������q� @B -C��6?0.1m     ��������q� ���� True     ��������q� ����  F     ��������q� ���� true     ��������q� ����  false     ��������               
                 q� ����     @�@1K      ��������q�  ����       ��������q�  ����       ��������q�  ����       ��������               
         ��              q�  ����        ��������              
                  q�  ����        ��������              
                                  
                 q�@ ����        ��������q�@ ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ���� true	     ��������q� ����  false
     ��������q� ���� true     ��������q� ����  false     ��������               
                 q� ����       5      ��������q� ����       5     ��������q� ����       5     ��������q� ����       5     ��������q� ����       ��������q� ����  	     ��������q� ����  
     ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ���� true     ��������q�@ ����       ��������q�@ ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����dec     ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ���� true     ��������q� ���� true     ��������q� ���� true     ��������q� ����  false     ��������q� ���� true     ��������q� ����  false      ��������q� ���� true!     ��������q� ����  false"     ��������               
                        q� ����       5      ��������q� ����       5     ��������q� ����       5     ��������q� ����       5     ��������q� ����       ��������q� ����  	     ��������q� ����  
     ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ���� true     ��������q�@ ����       ��������q�@ ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����dec     ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ���� true     ��������q� ���� true     ��������q� ���� true     ��������q� ����  false     ��������q� ���� true     ��������q� ����  false      ��������q� ���� true!     ��������q� ����  false"     ��������               
                 q� ����       5      ��������q� ����       5     ��������q� ����       5     ��������q� ����       5     ��������q� ����       ��������q� ����  	     ��������q� ����  
     ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ���� true     ��������q�@ ����       ��������q�@ ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����dec     ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ���� true     ��������q� ���� true     ��������q� ���� true     ��������q� ����  false     ��������q� ���� true     ��������q� ����  false      ��������q� ���� true!     ��������q� ����  false"     ��������               
                 q� ����       5      ��������q� ����       5     ��������q� ����       5     ��������q� ����       5     ��������q� ����       ��������q� ����  	     ��������q� ����  
     ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ���� true     ��������q�@ ����       ��������q�@ ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����dec     ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ���� true     ��������q� ���� true     ��������q� ���� true     ��������q� ����  false     ��������q� ���� true     ��������q� ����  false      ��������q� ���� true!     ��������q� ����  false"     ��������               
                 q�@ ����        ��������q�@ ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����decade     ��������q� ���� true     ��������q� ���� true     ��������q� ���� true     ��������q� ����  false     ��������               
                 q� ����        ��������q� ����       ��������q�@ ����       ��������q�  ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������q� ����       ��������               
                        q� ����dec     ��������q� ����     @�@1k     ��������q� ����    ��.A1meg     ��������q� ����       20     ��������q� ����        0     ��������q� ����        0     ��������q� ���� true	     ��������q� ���� true
     ��������q� ����      I@50     ��������q� ���� true     ��������q� ����  false     ��������               
                         / q� ���� x'     ��������q�     �-���q=1E-12     ��������q� @B -C��6?1E-4     ��������q� ���� x     ��������q� ���� x     ��������q� ���� x     ��������q� ���� x     ��������q� ���� x     ��������q� ���� x     ��������q� ���� x	     ��������q� ���� x!     ��������q� ����    �  500
     ��������q� ���� x     ��������q� ����    �  500     ��������q� ���� x$     ��������q� ���� x$     ��������q� ���� x%     ��������q� ���� x"     ��������q�  ���� x*     ��������q� ���� x     ��������q� ���� x     ��������q� ���� x     ��������q� ���� x&     ��������q� ���� x     ��������q� ���� x     ��������q� ���� x     ��������q� ���� x+     ��������q� ���� x,     ��������q� ���� x-     ��������q� ���� xg     ��������q� ���� xf     ��������q� ���� xd     ��������q� ���� xe     ��������q� ���� xh     ��������q� ���� xj     ��������q� ���� xi     ��������q� ���� xk     ��������q� ����    e��A1Gl     ��������q�             0�     ��������q� ����      @5�     ��������q� ����      @2.5�     ��������q� ����      �?.5�     ��������q� ����      @4.5�     ��������q� 
   ��&�.>1n�     ��������q� 
   ��&�.>1n�     ��������q� 
   ��&�.>1n�     ��������q� 
   ��&�.>1n�     ��������                 ���  CMacroBehavior      123 � � � buz-11buz-11 #               � � � MOSFETs   Siemens	   X5X5          ��*******
*n-mosfet*50v 30a 40mohm*add_in_line
.subckt buz-11 1  2  3
*pin order     g s d
ls 5 2 7n
ld 86 3 5n
rg 4 11 5.5m
rs 5 76 22m
d11 76 86 drev
.model drev d cjo=1.5n rs=20m tt=4.2n is=300p bv=50
m11 95 11 76 76 mbuz
.model mbuz nmos vto=3.315 kp=24.41
m2 11 95 8 8 msw
.model msw nmos vto=0.001 kp=5
m3 95 11 8 8 msw
cox 11 8 3n
dgd 8 95 dcgd
.model dcgd d cjo=1.03n m=0.537 vj=1.135
cgs 76 11 1.22n
m347 86 95 95 95 mvrd
.model mvrd nmos vto=-15.6 kp=10.5
lg 4 1 7n
.ends
                 Ariald     ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j                   ����            ��d               ��  TSignal                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                      	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CDCsweep       
 123456789:               
                       ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                       	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CACsweep        KLMNOPQR               
                       ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                      	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  �� 
 CTranSweep       ijklmnop               
                       ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                       	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CACdisto        defgh               
                           ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                       	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  c�        q� ����        ��������q� ����       ��������q� ����       ��������q� ����dec     ��������q� ����       ��������               
                           ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                       	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  c�        q� ����        ��������q� ����       ��������q� ����       ��������q� ����dec     ��������q� ����       ��������               
                           ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                       	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  c�        q� ����        ��������q� ����       ��������q� ����       ��������q� ����dec     ��������q� ����       ��������               
                           ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                       	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  c�        q� ����        ��������q� ����       ��������q� ����       ��������q� ����dec     ��������q� ����       ��������               
                           ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                       	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  c�        q� ����        ��������q� ����       ��������q� ����       ��������q� ����dec     ��������q� ����       ��������               
                       	    ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                      	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CACnoise        STUVWXYZ               
                    
    ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                      	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��         q�  ����        ��������q�  ����       ��������q�  ����       ��������q� ����dec     ��������q� ����       ��������q� ����       ��������q� ����  	     ��������q� ����  
     ��������              
                        ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                      	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CFourier        qrst               
         ��                   ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                      	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CACpz        	 [\]^_`abc               
                       ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                      	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CDCtf         ;<=>?               
                       ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                      	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CDCsens         @ABCDEFGHIJ               
                       ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                       	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j                  ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                      	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CShow         u              
                       ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                      	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CShowmod         v              
                       ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                      	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  �� 
 CLinearize        q�  ����        ��������               
                       ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                      	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CParamTranSweep        wxyz{|}~����               
                       ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                      	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  O              ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                       	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CParamACSweep        ������������                
                       ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                      	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CMonteCarlo_op        ����������������������������               
                              ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                      	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CMonteCarlo_dc        ����������������������������               
                       ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                       	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CMonteCarlo_ac        ����������������������������               
                       ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                      	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CMonteCarlo_tran        ����������������������������               
                       ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                       	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CACsens        	
               
                              ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                       	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CNetworkAnalysis                       
                       ����            P               H�                        v(1)       ����                  H�                       v(2)       ����                  H�                       v(3)       ����                  H�                       i(v1)       ����                  H�                       	v(i1_vrl)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j                  ����            P                 >           ��   CDigSimResTemplate                ���       ����  ����:�0�yU>20.00n���   ����                       Arial����                       Arial����                       Arial  �   �  �                                ����  ���� ������       ����  ���� ������                 �               ����  �����       200������         0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial      �       �         �     �   �  �  Circuit1                  ����  ��    ��������                        A                                                                                   A                             A                             A                    �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D �i�                T 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                      �  �                ր         �  @                  ���                                                  �  @  &�     <   �  <     ��                                                        &�     |   �  |     ��                                                        &�     �   �  �     ��                                                        &�     �   �  �     ��                                                        k� �      �  4     ��                                                      �      �  4   �      �  4   [title]                                       k� �   D   �  t     ��                                                      �   D   �  t   �   D   �  t   [description]                                       k� `   �   h  �     ��                                                      `   �   h  �   `   �   h  �   [id]                                       k� �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       k�      �   8    ��        	                                                   �   8       �   8  Date :       �    H  �                  k� �     �  4   	 ��        
                                              �     �  4  �     �  4  [date]                                       k�       t   8    
 ��                                                            t   8         t   8   Title :       �       �                  k�    L   �   x     ��                                                         L   �   x      L   �   x   Description :       �  �  �  �                  k�    �   �   �     ��                                                         �   �   �      �   �   �   ID :       �  �  �  P                  k�    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �  \  8                     ./012345689:;<          7     	title box    Analog Misc      �?    9 
 ԁ     q�  ����        ��������q�  ����       ��������q�  ����       ��������q�  ����       ��������q�  ����       ��������        9                                      ����؁�� ����     ځ            title                ځ            description               ځ            id               ځ            designer               ځ            date                           ����            `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                                                                                            2         �  �              � � �                   ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                        �   ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    
cgs 76         47 80moh5.6 B<
G7   mvrd nmodel 5   �@
G�
     H�                      TIME� # ) time                      H�                        i(v1)� < � i(v1)    TIME                 H�                        v(3)      v(3)    TIME                 H�                      	i(va_ix1)�   � 	i(va_ix1)    TIME                 H�    (v(3)-v(6))                  v(IVm1)� �   v(IVm1)    TIME                 H�                        v(6)      v(6)    TIME                           2         �  �           Time  � � �             ���
    ����                       Arial����                       Arial                              ����  �����z�`?2.035181e-003��G�6      ����  �����z�`?2.035181e-003��G�6      ����  ����1��{��%�-1.075922e+001������      ����  ����1��{��%�-1.075922e+001������                                                                       �                      �                                                                                                                                                                                                                                                                                                                                                                                                                              �                      �                                                                                                              �                      �                                                                                                              �                      �                              1m  0                            100   100                                                             1m  0                            100   100                                1m  0                            100   100                                1m  0                            100   100                                                 
                 1m  0                            100   100                                ��   CMiniPartPin    ����V+V+     PWR+V+g      Q�   ����V-V-     PWR-V-h     voltage_sourcevoltage_source                          Q�    ����Gate1     PASGateu      Q�   ����Source2     PASSourcew     Q�   ����Drain3     PASDrainv     BUZ11BUZ11                                  Q�    ����11     PAS1�      Q�   ����22     PAS2�     BatteryBattery                          Q�    ����R+R+     PASR+      Q�   ����R-R-     PASR-     RR                          Q�    ����GndGnd     GNDGnd}      GndGnd                  Q�    ����M+M+     PASM+i  4  Q�   ����M-M-     PASM-j  4  	voltmeter	voltmeter                          Q�    ����M+M+     PASM+2      Q�   ����M-M-     PASM-3     Ammeter2Ammeter2                          Q�    ����Gate1     PASGateu      Q�   ����Source2     PASSourcew     Q�   ����Drain3     PASDrainv     BUZ11BUZ11                                  Q�    ����V+V+     PWR+V+g      Q�   ����V-V-     PWR-V-h     voltage_sourcevoltage_source                          Q�    ����Gate1     PASGateu      Q�   ����Source2     PASSourcew     Q�   ����Drain3     PASDrainv     BUZ11BUZ11                                  Q�    ����V+V+     PWR+V+g      Q�   ����V-V-     PWR-V-h     voltage_sourcevoltage_source                          Q�    ����Gate1     PASGateu      Q�   ����Source2     PASSourcew     Q�   ����Drain3     PASDrainv     BUZ11BUZ11                                  Q�    ����V+V+     PWR+V+g      Q�   ����V-V-     PWR-V-h     voltage_sourcevoltage_source                                                                                                                                                
m1     8 8 mm l=100u w                        used                                                                                                                                                                                            (f    x=f � �'f                           �(f                            ,�e    �f � ��e                           ��e                                     �  � ���� �                         .I                                                                                                       
m1     8 8 mm l=100u w                        used                            tin    SSAGE: abortin
                        AGE:                            5011    53E-002
JV1.I y                        x��                              �@    �'@
G5   �@
G3                         ATAB                              �@    ��@
G5   �@
G3                         ATAB                            
>EN    A
>DATAB 5.01488                        A_IX    2 2 2 2 d                                                           