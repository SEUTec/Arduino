    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz        ��  CPart           �   �          �   �              Battery��  CIntPin    ��  CWire     �        �       �   �  �       �   �  �               resistor_generic �   �    �    
    �       �   �  �       �   �  �               resistor_generic �   �    �       �       _      �      _      �              capacitor_generic �   �     �         �           �   �           �   �               Gnd ��  CExtPin    ��  CVertex      �
   ��  CSegment/   �%      �	                  �5   �&   �  �
   �   �5   �  @                            �#    �>   @  �
   �6   �   @   
   "          !       �   ! �+   �
  �
   �"   �8   �
   
   &          %     �!   % �4   �  �
   �.   �   �  �   *     	    )     (          $                               `       Gnd}   �  �
          gnd1     ��   CPin                    ��                                                               Gnd��  TLine                   ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        .�         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        .�    ,   4   ,     ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        .�    8   (   8     ��    p�Z         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         - / 0 2   1      Ground    
Ground DINMiscellaneous      �?       ��   CGroundBehavior       Gnd ��   CBehPin     Gnd        ����Gnd����                        ��gndgnd                 6 Analog Meters   Generic   gnd1gnd1          ����  gnd ��   CPartPin    ����GndGnd      GNDAGnd    ����SourcesGroundGeneric              0 �         �       _   @  �      _   @  �              Ammeter29 �   �    �   <    3 ;  5�    2      ����2����                        ��5� �  M-      R  M-����                        �� 3  : 3 �        `   �  M+    �   �$      @   �4   �          C        B              `   `   M-    �  �        Isource    	 ,�                    ��                                                           �   M+,�                   ��                                                              M-.�     �       �     ��    ���                                                 .�     <             ��                                                        �� 
 TRectangle �����   @   <                  ����                                         ����<   @   �   .� ����x   ����L     ��    ���                                                 ��  TPolygon @�������@�������  ��          @ @                                           ��  TPoint����H    RGE.N�����T    �6�@N�����T       
@ @ ��  
 TTextField ����D   <   |     ��                                                      ����D   <   |   ����D   <   |   [value]       �  �  �  B	     D   �   |   R�    �����        ��                                                          �����         �����      	[refname]       �  �    h     �����      
 E F G H J S   K T M 	     Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       ��   CAmmeterBehavior     ��  CValue ?�]   @�p�? 9.00m      �������� M+M- 5� �  M+        R  M+����                        ��? AmmeterAmmeter   LD            Y ? Analog Meters   Generic   IsourceIsource          ����  VAm 7�    ����M+M+      PASAM+ 	X    7�   ����M-M-      PASAM-      Analog MetersAmmeter-verticalGeneric              0 �       �       _   �  �      _   �  �              
Voltmeter2�        ] 4 \ �    �=   �  �   �   �'   �  �   a �   b �A      �   �   �*      �   �'   �-      �   g �   h �0   �
  �   i                 f     e �   f �2   �  �   �,   l �   �  �   m    	        k             d     c �   �#   �  �   o         d                     `                `   `   M+    �      `   �  M-       `          Vsource    
 ,�                    ��                                                               M+,�                   ��                                                          �   M-.�     �       �     ��    ���                                                 .�             <     ��    �3V                                                .�    $      4     ��    ���                                                 .�    ,      ,     ��    (�K                                                .�    �      �     ��               	FIXED_ROT                                        I�     <   �   �                  ����                                             <   �   �   R�    D   �   x     ��                                                         D   �   x      D   �   x   [value]       ,  ,  $  �     D   �   x   R� 8      �   0    	 ��        	                                               8      �   0   8      �   0   	[refname]       �  �  H  $  8      �   0    r s v w x y z     {       u   t 
     Voltemeter-Vert    Voltemeter-Vert_smallMiscellaneous      �?       ��   CVoltmeterBehavior     W� ����      (@12.00      �������� M+M- 5� 4  M+        �  M+����                        ��5� 4  M-      �  M-����                        ��	voltmeter	voltmeter   X             � Analog Meters   Generic   VsourceVsource          ����  IVm 7�    ����M+M+      PASAM+ 
     7�   ����M-M-      PASAM-       Analog MetersVoltmeter-verticalGeneric              0  �        �       _      �      _      �              capacitor_generic�    �    �   �   �	       �      �      �      �              ua555�    �    � �   �   �       S   �  ,      S   �  ,              Ammeter�        � 4 � �    p        �   M+    �   �"   �  �   �   � �?   �  �   �    	                  �  �   M-    �  �          I555    	 ,�                   ��                                                           @   M+,�                   ��                                                      �   @   M-.� �   @   �   @     ��    ���                                                 .�     @       @     ��                                                        .� 4   X   `   X     ��    ���                                                 I�        �   d                   ����                                                �   d   L� ����������������  ��          @ @                                           N�d   X    �z�hN�X   P    C�mN�X   `    A��@ @ R� $   $   �   L     ��                                                      $   $   �   L   $   $   �   L   [value]       L  L  |  �  $   $   �   L   R�     �����        ��                                                           �����          �����      	[refname]       @  �     \      �����       �   � � �   �   � � �   � 	     Ammeter    Ammeter_smallMiscellaneous      �?       U�     W� ׀.   ��́? 8.69m      �������� M+M- 5� �  M+        R  M+����                        ��5� �  M-      R  M-����                        ��AmmeterAmmeter   W            � � Analog Meters   Generic   I555I555          ����  VAm 7�    ����M+M+      PASAM+h?W    7�   ����M-M-      PASAM-�YY   Analog MetersAmmeterGeneric              7  5�     vcc����    ����vcc����                        ���  7   � 7 �      � 5 � �      � 5 �      � 4 �   
   � 6 �   �    �    �    �   /   �      �   /   �      �               Marker� �    �<   �  `   �-   �   �  `   �    	    �                `      M     `  @         Vout     ,�                   ��                                                           `   M.� 0   `       `     ��    ���                                                 L� �����  �����     ��                                                         N�P   `    pQN�@   P       N�0   `        N�@   p            R� `   P      t     ��                                                       `   P      t   `   P      t   	[refname]       �  0  X  �        �   ,    �   � � �  �  Marker     Miscellaneous      �?    +   ��   CMarkerBehavior     W�             0.0      �������� M ��  	 TModelPin ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               � Analog MiscV   Generic   VoutVout          ����               Vout  v(Vout)  N 7�    ����MM       A    ����RootmarkerGeneric              Vout �  5�    out����   ����out����                        ���  Vout  � Vout �       � 0 �    �           VCC:  �   �3   �      �)   �.   @      � �7   �;   @  `   �3   � �	   �
  `   � �2   � �:   @  `   �                    �     �     �(   � �@   @  �   �+   � �   �  �   �    	        � �&   � �    @  @   �                        �        	          �  	THRESHOLD;  �   �   �  `   �*   �1   �
  `   � �    � �7   �
  @   �                �        	          �  Control<  �   �       @  TRIGGER=  �   n         RESET>  �   �   �      �0   � �6   `      � �   �9   `  `   �1   �
   `  `   �         �     �$   �,   `  �   �%   �/   `  �   �        �     �     �     �     �                	         �  	DISCHARGE?  �   �      �  OUTPUT@  �   +      @  GROUNDA   �  �          U1     ,�                    ��                                                           `   VCC,�                   ��                                                          �   	THRESHOLD,�                   ��                                                          �   Control,�                   ��                                                          �   TRIGGER,�                   ��                                                         `   RESET,�                   ��                                                         �   	DISCHARGE,�                   ��                                                         �   OUTPUT,�                   ��                                                         �   GROUND.�     `       `    	 ��                                                        .�     �       �    
 ��        	                                                .�     �       �     ��        
                                                .�     �       �     ��                                                        .� �   `      `     ��                                                        .� �   �      �     ��     ��                                                .� �   �      �     ��                                                        .� �   �      �     ��     �                                                 I�     @   �   �                  ����                                             @   �   �   R� (   P   p   p     ��                                                      (   P   p   p   (   P   p   p   vcc         p  �  �  (   P   p   p   R� (   p   p   �     ��                                                      (   p   p   �   (   p   p   �   thr         �  x  R  (   p   p   �   R� (   �   p   �     ��                                                      (   �   p   �   (   �   p   �   cont         0  �  �  (   �   p   �   R� (   �   p   �     ��                                                      (   �   p   �   (   �   p   �   trIg         �  �    (   �   p   �   R� �   P   �   p     ��                                                      �   P   �   p   �   P   �   p   reset       8  p  �  �  �   P   �   p   R� �   p   �   �     ��                                                      �   p   �   �   �   p   �   �   dischg       8  �  (  R  �   p   �   �   R� �   �   �   �     ��                                                      �   �   �   �   �   �   �   �   out       8  0  �  �  �   �   �   �   R� �   �   �   �     ��                                                      �   �   �   �   �   �   �   �   gnd       8  �  �    �   �   �   �   R�     �����        ��                                                           �����          �����      	[devname]        ����������������    �����      R�        �   <     ��                                                              �   <          �   <   	[refname]          �  �  h         �   <    � � � � � � � � �   � � � � � � � � � � � � �  �      lm555     Miscellaneous      �?   #    U 7�    ����VCCvcc      PASAVCC    ����7�   ����	THRESHOLDthr      PASA	THRESHOLD    ����7�   ����Controlctrl      PASAControl    ����7�   ����TRIGGERtrg      PASATRIGGER��S����7�   ����RESETrst      PASARESET�<
����7�   ����	DISCHARGEdis      PASA	DISCHARGE    ����7�   ����OUTPUTout      PASAOUTPUT�eR����7�   ����GROUNDground      PASAGROUNDDANA����Timer	555 timerNational Semiconductor              8 �  5�    ctrl����   ����ctrl����                        ��5�     C+        ����C+����                        �� 8  � 8 � �    '       �  C-�P�   �        �   C+ �  �
  �         Cc     ,�                   ��                                                           �   C-,�                   ��                                                          @   C+.�     @       �      ��                                                        .�     �   �����     ��                                                        .�     �   �����     ��                                                        .�     �       �     ��                                                        R� 0   t   �   �     ��                                                       0   t   �   �   0   t   �   �   [capacitance]         �  �  r	      `   �   �   R� 0   @   �   d     ��                                                       0   @   �   d   0   @   �   d   	[refname]         @  �  �          �   $               �  	Capacitor     Miscellaneous      �?       ��  CCapacitorBehavior     W� '  ��&�.>1n      ��������W� ���� x     ��������W� ����       ��������W� ����       �������� C+C- 5�    C-      ����C-����                        �� 	capacitor   i            Passive   Generic   CcCc          ����  C 7�    ����C+C+      PASAC+   �����7�   ����C-C-      PASAC-    ����Passive Generic              0 �  6 5�    C-      ����C-����                        ��5�    ground����   ����GROUND����                        ��� Y   0     0 �    #       �  C-�  �   �        �   C+�   @  �         C1     ,�                   ��                                                           �   C-,�                   ��                                                          @   C+.�     @       �      ��    
*                                                 .�     �   �����     ��     gro                                                .�     �   �����     ��     
q                                                .�     �       �     ��    jt_n                                                R� 0   t   �   �     ��                                                       0   t   �   �   0   t   �   �   [capacitance]       �  �  x	  r	      `   �   �   R� 0   @   �   d     ��                                                       0   @   �   d   0   @   �   d   	[refname]       �  @  P	  �          �   $    '()*+    ,      %& �  	Capacitor     Miscellaneous      �?       �     W� '  +�|�;i>47n      ��������W� ���� x     ��������W� ����       ��������W� ����       �������� C+C- 5�     C+        ����C+����                        ��! 	capacitor   i            2!Passive   Generic   C1C1          ����  C 7�    ����C+C+      PASAC+��X����7�   ����C-C-      PASAC-    ����Passive Generic              5 � �   25�    R-      ����R-����                        ��5�    thr����   ����thr����                        ��5�    trg����   ����trg����                        �� 5   5 �    �    �  �   R+  �   �       �   R-   �
  �         R2     ,�                    ��                                                       �   @   R+,�                   ��                                                          @   R-.�    @   $   0     ��    �                                                 .� 0   P   $   0     ��                                                       .� 0   P   <   0     ��    ��K                                                .� H   P   <   0     ��                                                       .� H   P   T   0     ��                                                        .� `   P   h   @     ��    (�K                                                .� �   @   h   @     ��                                                       .� `   P   T   0    	 ��        	                                                .�    @       @    
 ��        
                                                R�     `   �   �     ��                                                           `   �   �       `   �   �   [resistance]       �
  �  �  V      `   �   �   R�         t   $     ��                                                               t   $           t   $   	[refname]       �
  �  `  @          t   $    :;<=>?@ABCDEF   resistor    resistor DINMiscellaneous      �?       ��  CResistorBehavior     W� ����     ��@10k      ��������W� ���� 27     ��������W� ����       ��������W� ����       �������� R+R- 5�     R+        ����R+����                        ��5 resistor   i            M5Passive   Generic   R2R2          ����    R 7�    ����R+R+      PASAR+DATA����7�   ����R-R-      PASAR-G3 ����Passive Generic              6 	 �  M5�    dis����   ����dis����                        ��5� �,  R-      
  R-����                        �� 6   6 �    j        �   R+    �   �   �  �   R-    �
             R1     ,�                    ��                                                           @   R+,�                   ��                                                      �   @   R-.� d   @   \   P     ��    ���                                                 .� P   0   \   P     ��                                                        .� P   0   D   P     ��    ���                                                 .� 8   0   D   P     ��    (�K                                                .� 8   0   ,   P     ��                                                       .�     0      @     ��    ��K                                                .�     @      @     ��                                                       .�     0   ,   P    	 ��        	                                                .� d   @   �   @    
 ��        
                                                R�     `   �   �     ��                                                           `   �   �       `   �   �   [resistance]       �
  @  �  �      `   �   �   R�         t   $     ��                                                               t   $           t   $   	[refname]       �
     `  �          t   $    TUVWXYZ[\]^_`     resistor    resistor DINMiscellaneous      �?       G�     W� ����     \�@4.7k      ��������W� ���� 27     ��������W� ����       ��������W� ����       �������� R+R- 5� �,  R+        
  R+����                        ��Q resistor   S           fQPassive   Generic   R1R1          ����    R 7�    ����R+R+      PASAR+   �    7�   ����R-R-      PASAR-       Passive Generic              4 � ^ �  5�     1       ����1����                        ��5�    rst����   ����rst����                        ���  f 4    4 = �    d    `       1�  �   D   `   �  2�   �  �          X1     ,�                    ��                                                               1,�                   ��                                                          �   2.�             $     ��    ��)                                                .�     \       �     ��                                                        .�    8   0   8    	 ��    ��)                                                .�     H   @   H     ��    p�Z                                                .�     $   @   $     ��                                                       .�    \   0   \     ��    D�Z                                                .�               ���                                                      .�               ���   �Z	                                                R� `          $    
 ��        
                                               `          $   `          $   	[devname]        ����������������`          $   R� `   $      H     ��                                                       `   $      H   `   $      H   	[refname]       �    P  �  `   $      H    mnopstuv    wx    r  q     Battery     Miscellaneous      �?    9 
 ��  CParamSubBehavior     W� ����      (@12      �������� 12 i> BatteryBattery
 9 i             i> Sources   Generic   X1X1          ������   CParamSubModelType��    BATTERY2.SUBCKT Xbattery 1 2
V1 1 2 DC {voltage}
.ENDS
   ��  	 CParmDefn    1battery voltage   ParamSubvoltageV                X 7�    ����11      PASA1�Y����7�   ����22      PASA2�1b����SourcesBatteryGeneric                       �   � ] :  � �     �  <  
 � � 8 " 8                                             � o  $ a e c k i � � ( &   � � � g � � � � m � *  � � � � C  " � B * B �       #        � � �               D             + �   n � �     � p B   b     f % � h � � j � l � )  � � ' � � � � ` ! � � d                    
 W�@ ����        ��������W�             0     ��������W� ����      @5     ��������W�  ʚ;�������?.1     ��������W�@ ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ���� true
     ��������W� ����  false     ��������               
                  W� ����        ��������W� ����       ��������W�  ����       ��������W�@ ����       ��������W�@ ����       ��������               
                  W� ����        ��������W� ����       ��������W�@ ����       ��������W�  ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������               
                 W� ����dec     ��������W� ����     @�@1k     ��������W� ����    ��.A1meg     ��������W� ����       20     ��������W� ���� true     ��������W� ���� true     ��������W� ���� true	     ��������W� ����  false
     ��������               
                 W�  ����        ��������W�  ����       ��������W�  ����       ��������W� ����dec     ��������W� ����       ��������W� ����       ��������W� ����  	     ��������W� ����  
     ��������               
                  	 W� ����        ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������               
                 W� ����        ��������W� ����       ��������W� ����       ��������W� ����dec     ��������W� ����       ��������               
                    W�             0      ��������W� ����~j�t�h?3m     ��������W� �� �h㈵��>10u     ��������W� �� �h㈵��>10u     ��������W� ���� True     ��������W� ����  F     ��������W� ���� true     ��������W� ����  false     ��������               
                 W� ����     @�@1K      ��������W�  ����       ��������W�  ����       ��������W�  ����       ��������               
         ��              W�  ����        ��������              
                  W�  ����        ��������              
                                  
                 W�@ ����        ��������W�@ ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ���� true	     ��������W� ����  false
     ��������W� ���� true     ��������W� ����  false     ��������               
                 W� ����       5      ��������W� ����       5     ��������W� ����       5     ��������W� ����       5     ��������W� ����       ��������W� ����  	     ��������W� ����  
     ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ���� true     ��������W�@ ����       ��������W�@ ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����dec     ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ���� true     ��������W� ���� true     ��������W� ���� true     ��������W� ����  false     ��������W� ���� true     ��������W� ����  false      ��������W� ���� true!     ��������W� ����  false"     ��������               
                        W� ����       5      ��������W� ����       5     ��������W� ����       5     ��������W� ����       5     ��������W� ����       ��������W� ����  	     ��������W� ����  
     ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ���� true     ��������W�@ ����       ��������W�@ ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����dec     ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ���� true     ��������W� ���� true     ��������W� ���� true     ��������W� ����  false     ��������W� ���� true     ��������W� ����  false      ��������W� ���� true!     ��������W� ����  false"     ��������               
                 W� ����       5      ��������W� ����       5     ��������W� ����       5     ��������W� ����       5     ��������W� ����       ��������W� ����  	     ��������W� ����  
     ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ���� true     ��������W�@ ����       ��������W�@ ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����dec     ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ���� true     ��������W� ���� true     ��������W� ���� true     ��������W� ����  false     ��������W� ���� true     ��������W� ����  false      ��������W� ���� true!     ��������W� ����  false"     ��������               
                 W� ����       5      ��������W� ����       5     ��������W� ����       5     ��������W� ����       5     ��������W� ����       ��������W� ����  	     ��������W� ����  
     ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ���� true     ��������W�@ ����       ��������W�@ ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����dec     ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ���� true     ��������W� ���� true     ��������W� ���� true     ��������W� ����  false     ��������W� ���� true     ��������W� ����  false      ��������W� ���� true!     ��������W� ����  false"     ��������               
                 W�@ ����        ��������W�@ ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����decade     ��������W� ���� true     ��������W� ���� true     ��������W� ���� true     ��������W� ����  false     ��������               
                 W� ����        ��������W� ����       ��������W�@ ����       ��������W�  ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������W� ����       ��������               
                        W� ����dec     ��������W� ����     @�@1k     ��������W� ����    ��.A1meg     ��������W� ����       20     ��������W� ����        0     ��������W� ����        0     ��������W� ���� true	     ��������W� ���� true
     ��������W� ����      I@50     ��������W� ���� true     ��������W� ����  false     ��������               
                         / W� ���� x'     ��������W�     �-���q=1E-12     ��������W� @B -C��6?1E-4     ��������W� ���� x     ��������W� ���� x     ��������W� ���� x     ��������W� ���� x     ��������W� ���� x     ��������W� ���� x     ��������W� ���� x	     ��������W� ���� x!     ��������W� ����    �  500
     ��������W� ���� x     ��������W� ����    �  500     ��������W� ���� x$     ��������W� ���� x$     ��������W� ���� x%     ��������W� ���� x"     ��������W�  ���� x*     ��������W� ���� x     ��������W� ���� x     ��������W� ���� x     ��������W� ���� x&     ��������W� ���� x     ��������W� ���� x     ��������W� ���� x     ��������W� ���� x+     ��������W� ���� x,     ��������W� ���� x-     ��������W� ���� xg     ��������W� ���� xf     ��������W� ���� xd     ��������W� ���� xe     ��������W� ���� xh     ��������W� ���� xj     ��������W� ���� xi     ��������W� ���� xk     ��������W� ����    e��A1Gl     ��������W�             0�     ��������W� ����      @5�     ��������W� ����      @2.5�     ��������W� ����      �?.5�     ��������W� ����      @4.5�     ��������W� 
   ��&�.>1n�     ��������W� 
   ��&�.>1n�     ��������W� 
   ��&�.>1n�     ��������W� 
   ��&�.>1n�     ��������                 z��  CMacroBehavior      vccthrctrltrgrstdisoutground � 67jP� "ua555ua555 # u             � 67jP� "Timer�   Generic   U1U1          ��************************
* B2 Spice Subcircuit
************************
* Pin #		Pin Name
* vcc		vcc
* thr		thr
* ctrl		ctrl
* trg		trg
* rst		rst
* dis		dis
* out		out
* GROUND		GROUND
.Subckt ua555 vcc thr ctrl trg rst dis out GROUND 


***** main circuit
R1 vcc  9  4.7K 
R2 vcc  3  830 
R3 vcc  8  4.7k 
R4 vcc  10  1K 
R5 vcc  ctrl  5K 
R7 17  0  10K 
Q6 2  thr  5 bjt_npn_generic 
Q2 25  2  3 bjt_pnp_generic 
Q3_ 0  6  3 bjt_pnp_generic 
Q1 2  2  9 bjt_pnp_generic 
Q7 2  5  17 bjt_npn_generic 
Q8 6  4  17 bjt_npn_generic 
Q9 6  ctrl  4 bjt_npn_generic 
Q4 6  6  8 bjt_pnp_generic 
Q5 12  20  10 bjt_pnp_generic 
Q17_ 15  rst  31 bjt_pnp_generic 
Q16 dis  15  0 bjt_npn_generic 
R14_ 15  16  100 
Q14_ 0  trg  11 bjt_pnp_generic 
Q12_ 22  11  12 bjt_pnp_generic 
Q13_ 14  13  12 bjt_pnp_generic 
Q15_ 14  18  13 bjt_pnp_generic 
R8_ 22  0  100K 
R0 ctrl  18  5K 
R10 18  0  5K 
Q21_ 25  22  0 bjt_npn_generic 
Q20_ 24  25  0 bjt_npn_generic 
Q22_ 27  24  0 bjt_npn_generic 
Q24_ 29  27  16 bjt_npn_generic 
Q25_ out  26  0 bjt_npn_generic 
Q23_ vcc  29  28 bjt_npn_generic 
Q26 vcc  28  out bjt_npn_generic 
Q19 20  20  vcc bjt_pnp_generic 
R11_ 20  31  5K 
D1 31  24 diode 
R12_ 25  27  4.7K 
R15_ 16  26  220 
R16_ 16  0  4.7K 
D2 out  29 diode 
R6_ vcc  29  6.8K 
R17_ 28  out  3.9K 
R9_ 14  0  100K 
Q18 27  20  vcc bjt_pnp_generic 

.model bjt_npn_generic npn  is = 5f   bf = 100    nf = 1   vaf = 160   ikf = 30m   ise = 4p  
+ ne = 2   br = 4   nr = 1   var = 16   ikr = 45m  
+ rb = 4   re = 1.0   rc = .4   cje = 12.4p   vje = 1.1  
+ mje = .5   tf = 250p   cjc = 4p   vjc = .3   mjc = .3  
+ tr = 1n  

.model bjt_pnp_generic pnp  is = 1.0e-14   bf = 20    vaf = 50   ne = 2   br = .02   rb = 25  
+ rc = 4   cje = 12.4p   vje = 1.1   mje = .5   tf = 250p  
+ vjc = .3   mjc = .3   tr = 100n  

.model diode D  is = 1.0E-14   rs = 40   cjo = 1p  

.ends                 Ariald     �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j                   ����            ��W               ��  TSignal                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��  CDCsweep       
 ����������               
                       ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��  CACsweep        ��������               
                       ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  �� 
 CTranSweep       ��������               
                       ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��  CACdisto        �����               
                           ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��        W� ����        ��������W� ����       ��������W� ����       ��������W� ����dec     ��������W� ����       ��������               
                           ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��        W� ����        ��������W� ����       ��������W� ����       ��������W� ����dec     ��������W� ����       ��������               
                           ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��        W� ����        ��������W� ����       ��������W� ����       ��������W� ����dec     ��������W� ����       ��������               
                           ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��        W� ����        ��������W� ����       ��������W� ����       ��������W� ����dec     ��������W� ����       ��������               
                           ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��        W� ����        ��������W� ����       ��������W� ����       ��������W� ����dec     ��������W� ����       ��������               
                       	    ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��  CACnoise        ��������               
                    
    ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��         W�  ����        ��������W�  ����       ��������W�  ����       ��������W� ����dec     ��������W� ����       ��������W� ����       ��������W� ����  	     ��������W� ����  
     ��������              
                        ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��  CFourier        ����               
         ��                   ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��  CACpz        	 ���������               
                       ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��  CDCtf         �����               
                       ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��  CDCsens         �����������               
                       ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j                  ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��  CShow         �              
                       ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��  CShowmod         �              
                       ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  �� 
 CLinearize        W�  ����        ��������               
                       ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��  CParamTranSweep        �������������               
                       ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  �              ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��  CParamACSweep        EFGHIJKLMNOPQ               
                       ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��  CMonteCarlo_op        ����������������������������               
                              ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��  CMonteCarlo_dc        ��������������� 	
               
                       ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��  CMonteCarlo_ac         !"#$%&'(               
                       ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��  CMonteCarlo_tran        )*+,-./0123456789:;<=>?@ABCD               
                       ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��  CACsens        RSTUVWXYZ[\               
                              ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j  ��  CNetworkAnalysis        ]^_`abcdefg               
                       ����            P               ��                        v(vout)       ����                  ��                       v(4)       ����                  ��                       v(3)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  �  �� �|p�|����m�|+j  �  �� �|p�|����m�|+j                  ����            P                 >           ��   CDigSimResTemplate                ���       ����  ����:�0�yU>20.00n���   ����                       Arial����                       Arial����                       Arial  �   �  �                                ����  ���� ������       ����  ���� ������                 �               ����  �����       200������         0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial      �       �         �     �   �  �  Circuit1                  ����  ��    ��������                                                                                                                                                                   �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            B  �                C K�� ��    E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                      �  �                I�         �  @                  ���                                                  �  @  .�     <   �  <     ��                                                        .�     |   �  |     ��                                                        .�     �   �  �     ��                                                        .�     �   �  �     ��                                                        R� �      �  4     ��                                                      �      �  4   �      �  4   [title]                                       R� �   D   �  t     ��                                                      �   D   �  t   �   D   �  t   [description]                                       R� `   �   h  �     ��                                                      `   �   h  �   `   �   h  �   [id]                                       R� �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       R�      �   8    ��        	                                                   �   8       �   8  Date :       �    H  �                  R� �     �  4   	 ��        
                                              �     �  4  �     �  4  [date]                                       R�       t   8    
 ��                                                            t   8         t   8   Title :       �       �                  R�    L   �   x     ��                                                         L   �   x      L   �   x   Description :       �  �  �  �                  R�    �   �   �     ��                                                         �   �   �      �   �   �   ID :       �  �  �  P                  R�    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �  \  8                     ��������������          �     	title box    Analog Misc      �?    9 
 y�     W�  ����        ��������W�  ����       ��������W�  ����       ��������W�  ����       ��������W�  ����       ��������        9                                      ����|��� ����     ~�            title                ~�            description               ~�            id               ~�            designer               ~�            date                           ����            `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                                                                                            2         �  �              � � �                   ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                            �   ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    
cgs 76         47 80moh5.6 >DATAB 2mvrd nmodel -003
MVIJV    	 ��                      TIME� # ) time                      ��                        v(3)      v(3)    TIME                 ��                        v(4)      v(4)    TIME                 ��                       v(vout)      v(vout)    TIME                 ��    v(4)                   
v(Vsource)� �   
v(Vsource)    TIME                 ��                       
i(isource)�   � 
i(isource)    TIME                 ��    v(vsource)*i(isource)                   Psource� �    ����TIME                 ��                       i(i555)� �   i(i555)    TIME                 ��    i(i555)*v(Vsource)                   P555� � �  ����TIME                           2         �  �           Time  � � �             548E    ����                       Arial����                       Arial                              ����  �����z�`?2.035181e-003��G�6      ����  �����z�`?2.035181e-003��G�6      ����  ����1��{��%�-1.075922e+001������      ����  ����1��{��%�-1.075922e+001������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           1m  0                            100   100                             100     100  1m0                   1m  0                            100   100                                1m  0                            100   100                                1m  0                            100   100                                                 
                 1m  0                            100   100                                ��   CMiniPartPin    ����11     PAS1�         ����22     PAS2�     BatteryBattery                              ����GndGnd     GNDGnd}      GndGnd                      ����C+C+     PASC+�         ����C-C-     PASC-�     capacitor_genericcapacitor_generic                              ����R+R+     PASR+         ����R-R-     PASR-     resistor_genericresistor_generic                              ����VCCvcc     PASVCC:         ����	THRESHOLDthr     PAS	THRESHOLD;        ����Controlctrl     PASControl<        ����TRIGGERtrg     PASTRIGGER=        ����RESETrst     PASRESET>        ����	DISCHARGEdis     PAS	DISCHARGE?        ����OUTPUTout     PASOUTPUT@        ����GROUNDground     PASGROUNDA     ua555ua555                                                                              ����M+M+     PASM+0  �     ����M-M-     PASM-1  �  AmmeterAmmeter                              ����M+M+     PASM+k  4     ����M-M-     PASM-l  4  
Voltmeter2
Voltmeter2                              ����M+M+     PASM+2  �     ����M-M-     PASM-3  �  Ammeter2Ammeter2                              ����R+R+     PASR+  �,     ����R-R-     PASR-  �,  resistor_genericresistor_generic                              ����C+C+     PASC+�         ����C-C-     PASC-�     capacitor_genericcapacitor_generic                              ����MM       ��������MarkerMarker                                                                                                                                                                                                                        ,�e    �f � ��e                           ��e                                        ! � ��t                                                        ����       �� <                                                                               �    �Q                        6                             ��Z    P�W��W��W8KX                        �_�                            �Y    P�W��W��W��W                        ��W                            �`?     � @�R �  �                          ��                                                                            ����                                     �  � ���� �                                                         B 2.    224912E-003
IOUT                           @    2 2 2 2 d                                                     