    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz    ��  CPart    �����   �  �  �����   �  �              voltage_source��  CIntPin    ��  CWire    �        �   /   �   �      /   �   �                  Marker ��  CExtPin    ��  CVertex   �
  @   ��  CSegment    �   �
   	                          `      M      
             VControl     ��   CPin                   ��                                                           `   M��  TLine     P       `     ��    ���                                                 ��  TPolygon     ����    ����   ��                                                         ��  TPoint    0    Amm�   @        �    P        �0   @    P�X    ��  
 TTextField       �   ,     ��                                                             �   ,         �   ,   	[refname]       8
  8  �  �        �   ,               Marker     Miscellaneous      �?    +   ��   CMarkerBehavior     ��  CValue             0.0      �������� M ��  	 TModelPin ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �         �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               " Analog MiscV   Generic   VControlVControl          ����               VControl  v(VControl)  N ��   CPartPin    ����MM       A  ������RootmarkerGeneric              VControl �        �   /   �   �      /   �   �                  Marker% 	�    �3   `  @   �   ( �2   `   	   )                       `      M                   VControl     �                   ��                                                           `   M�     P       `     ��    ���                                                 �     ����    ����   ��                                                         �    0        �   @    ����    P    H���0   @    ��    �       �   ,     ��                                                             �   ,         �   ,   	[refname]         8  �  �        �   ,    -   + 2 ,      Marker     Miscellaneous      �?    +   �     �             0.0      �������� M !� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      3   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               5 Analog MiscV   Generic   VControlVControl          ����               VControl  v(VControl)  N #�    ����MM       A Teu ����RootmarkerGeneric              VControl �        �	   /   �   �      /   �   �                  Marker7 	�    �4      �   �-   : �      �   ;                 	        `      M     �  �          VControl     �                   ��                                                           `   M�     P       `     ��    ���                                                 �     ����    ����   ��                                                         �    0      �   @      �    P        �0   @            �       �   ,     ��                                                             �   ,         �   ,   	[refname]       �  �  s  �        �   ,    ?   = D >      Marker     Miscellaneous      �?    +   �     �             0.0      �������� M !� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      E   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               G Analog MiscV   Generic   VControlVControl          ����               VControl  v(VControl)  N #�    ����MM       A     ����RootmarkerGeneric              VControl  �      �       �   �  �      �   �  �              vcswitch�    �     �    L     �           �   �           �   �               GndM 	�    �$   `  �   �!   �.   `  �
   Q         P     �    �8   �  �   �/   �   �  �
   U          T     S      P     �   P �/   �  �   �'   �   �  �
   Y          X     W �   X �5   �
  �   [ �   \ �,   @  �   ] �)   �   @  �
   _         ^              �&   �   �
  �
   a         \                                   `       Gnd}      �          gnd1     �                    ��                                                               Gnd�                   ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��    ���          AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��    ���          AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��    ��K         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         c d e g   f      Ground    
Ground DINMiscellaneous      �?       ��   CGroundBehavior       Gnd ��   CBehPin     Gnd        ����Gnd����                        ��gndgnd                 k Analog Meters   Generic   gnd1gnd1          ����  gnd #�    ����GndGnd      GNDAGnd    ����SourcesGroundGeneric              0 �   L    J 0 K �    L     �       _   @  �      _   @  �              Ammeter2n �   �    �   q   �           �   �          �   �              Battery�    �    �    u    �   /   �      �   /   �      �               Markerv 	�    �+   �  `   �   �   �      z         y     �   �&   �  @   �   �;   @  @   ~         }     �,   �9   �  @   �    
     }     |     y                `      M     `  @         VSource     �                   ��                                                           `   M� 0   `       `     ��    ���                                                 �     `       `      ��                                                         �P   `    �F��@   P    G8 ��0   `    .383�@   p    E.I     � `   P      t     ��                                                       `   P      t   `   P      t   	[refname]       �  0  	  �        �   ,    �   � � �  �  Marker     Miscellaneous      �?    +   �     �             0.0      �������� M !� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     u �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  + X5            � Analog MiscV   Generic   VSourceVSource          ����               VSource  
v(VSource)  N #�    ����MM       A I ������RootmarkerGeneric              VSource t �    u    �       �   �        �   �                Inductor� �   �    �   �   �       �   �  �      �   �  �              	voltmeter�    �    � �   �   �
       �   �        �   �                Inductor�    u    � VSource � 	�    �    �  �   L+K  	�   �1   �  @   �   �0   �  @   � �%   �"   �      �   � �%   �      �             �     �     �   � �*   �      �(   � �6   �      � �$   � �7   @      �                     �   � �   �  �   �             �             �        
          �   L-L   �  �         L2     �                    ��                                                       �   @   L+�                   ��                                                          @   L-��   TArc ,����  T����   
                                                               ,   8   T       ,   8   T       @   8   @           �� ,���p  T����   	                                                           8   ,   P   T   8   ,   P   T   8   @   P   @           �� ,���X  T���p                                                              P   ,   h   T   P   ,   h   T   P   @   h   @           �� ,���@  T���X                                                              h   ,   �   T   h   ,   �   T   h   @   �   @           � |   0   �   (     ��    t                                                � �   8   |   0     ��     "                                                 � �   0   |   0     ��                                                        � �   @   �   @     ��    ���	                                                �     @   ����@     ��    ����
                                                �     \   �   |     ��                                                           \   �   |       \   �   |   [Inductance]       �  �  2  "      \   �   |   �         �   $     ��                                                               �   $           �   $   	[refname]       �  �  2  +          �   $    � � �   �   �   �   � � �   �   �   �   �    Inductor     Miscellaneous      �?    
   ��  CInductorBehavior     � ��� {�G�zt?5m      ��������� ���� x     �������� L+L- j�     L+        ����L+����                        ��j�    L-      ����L-����                        �� Inductor  
 �           � � Passive   Generic   L2L2          ����  L #�    ����L+L+      PASAL+    ����#�   ����L-L-      PASAL-    ����PassiveInductorGeneric              3 �   �    �       _   �         _   �                 capacitor_generic�    �   � 4 � 	�    �       �   C-�  	�   �-   �	      �"   � �(   @      � �   �)   @  @   �   �:    
  @   �        �     �#   �!   @      �   �#   @      �        �     �     �     �     �     �   � �   @  �   �                               �  �   C+�   �  `         C1     �                   ��                                                           @   C-�                   ��                                                      �   @   C+� �   @   `   @      ��    ��                                                � `   `   `         ��                                                        � @   `   @         ��    ��                                                � @   @       @     ��    p�H                                                �     `   �   �     ��                                                           `   �   �       `   �   �   [capacitance]       �  �  �        `   �   �   �         �   $     ��                                                               �   $           �   $   	[refname]       �  `  i            �   $    � � � � �     �       � �    	Capacitor     Miscellaneous      �?       ��  CCapacitorBehavior     � '  -C��6?0.1m      ��������� ���� x     ��������� ����       ��������� ����       �������� C+C- j�     C+        ����C+����                        ��j�    C-      ����C-����                        �� 	capacitor   N           � � Passive   Generic   C1C1          ����  C #�    ����C+C+      PASAC+    ����#�   ����C-C-      PASAC-    ����Passive Generic              3 �    �    �       _   @  �      _   @  �              Ammeter2� �   �    � �    �    �       �   �         �   �                 1n4007� �   �    �   �   J 7 �  j�    2      ����2����                        ��j�   D-      (  D-����                        �� 7  � 7 	�    �   �      �   � �   �  `   �                              D+    	�   �   �  @   �   � �   �   	   �                         @  D-    �            D1     �                   ��                                                           `   D+�                   ��                                                          �   D-�     �       �      ��    ���                                                 �     �   �����     ��                                                        �     �   �����     ��    ���                                                 �     `       �     ��                                                       �    �       �     ��    ��K                                                �     �   �����     ��    ��K                                                �     �       �     ��                                                        � 0   `   �   �    	 ��        	                                               0   `   �   �   0   `   �   �   	[devname]        �������������������������      � 0   �   �   �    
 ��        
                                               0   �   �   �   0   �   �   �   	[refname]       0  �  �  g  ����   �   <    � � � � � � �                � �  �  diode     Miscellaneous      �?       ��  CDiodeBehavior     � ����        ��������� ���� 27     ��������� ����       ��������� ����       �������� D+D- j�   D+        (  D+����                        ��� d1n4007d1n4007    �          � Diode   Generic   D1D1                D #�    ����D+D+      PASAA@�    #�   ����D-D-      PASAK�l   DiodeDiode	FairchildDO-41             9  j�    M-      ����M-����                        �� 9  � 9 	�    �    `   `   M+2  	�   �   `   �  M-3   @  �        IS1    	 �                    ��                                                               M+�                   ��                                                          �   M-�             <     ��     T                                                �     �       �     ��                                                        �� 
 TRectangle �����   @   <                  ����                                         ����<   @   �   � ����H   ����t     ��                                                        �  ������� �������  ��          @ @                                           �����x    ��b�����l    
>DA�����l    uT@ @ � ����D   <   |     ��                                                      ����D   <   |   ����D   <   |   [value]         L  =  �     D   �   |   � ��������B        ��                                                       ��������B      ��������B      	[refname]       �   b  f       �����      
   	   Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       ��   CAmmeterBehavior     � �w    @�%?160.35u      �������� M+M- j�     M+        ����M+����                        ��AmmeterAmmeter   V            Analog Meters   Generic   IS1IS1          ����  VAm #�    ����M+M+      PASAM+�������#�   ����M-M-      PASAM-������Analog MetersAmmeter-verticalGeneric              3  j�     M+        ����M+����                        ��� �  3   � 3 � 	�    �           M+i  	�   �   �     M-j   �              Vp    
 �                   ��                                                           `   M+�                   ��                                                      �   `   M-�     `       `     ��    ���                                                 � �   `   �   `     ��                                                       �    L      \     ��    ���                                                 �     T      T     ��    (�K                                                � �   X   �   X     ��               	FIXED_ROT                                        �     <   �   �                   ����                                             <   �   �   � (   D   �   x     ��                                                      (   D   �   x   (   D   �   x   [value]         �     Z  (   D   �   x   �        �   0    	 ��        	                                                      �   0          �   0   	[refname]          $   ~  �          �   0    +  $%&,(  )-*      '
     	voltmeter    voltmeter_smallMiscellaneous      �?       ��   CVoltmeterBehavior     � ����    �0�-16.01      �������� M+M- !j�    M-      ����M-����                        ��	voltmeter	voltmeter   �            !1Analog Meters   Generic   VpVp          ����  IVm #�    ����M+M+      PASAM+- � ����#�   ����M-M-      PASAM-NAL
����Analog Meters Generic              4 � � �    �    �       _   @  �      _   @  �              Ammeter24�   �	    6�    7  	 �       �   �         �   �                 1n40078�   �    �    ;   �       �   �  �      �   �  �              vcswitch<�   L    =0 �   L    =0 �      =VControl 	�    �   @   	   �   �   @  @   C       B               �      1S  	�   `   �   �  2T  	�   b       �  3U  	�             4V   �
  �       X4     �                    ��                                                       @   `   1�                   ��                                                      @   �   2�                   ��                                                          �   3�                   ��                                                          `   4�     �       `     ��    ��                                                �     �       �     ��                                                        �     �       �    
 ���   ��                                                � �����      �    	 ���   p�H                                                ��  TEllipse <   �   D   �                  ����                                         <   �   D   �   <   �   D   �   � �����      �               	   ����                                         �����      �   � @   �   @   �     ��       
                                                � 0   �   @   �     ��    D�H                                                � @   �   @   `     ��                                                       �    �   �����     ��  � �H        	FIXED_ROT                                        �    �   4   �     ��    .I                                                  � `   �   �   �     ��                                                       `   �   �   �   `   �   �   �   	[refname]       �  �	    G
      (   t   L   � `   `   �   �     ��                                                       `   `   �   �   `   `   �   �   	[devname]        ����������������       �   (    HIJKRSU      MV  WOXYTLN    Q �  vcswitch     Miscellaneous      �?   9 
 ��  CParamSubBehavior    � ����      @3      ��������� ����      @3     ��������� ����      �?0.5     ��������� ����    ��.A1meg     �������� 1234 j�     1       ����1����                        ��j�    2      ����2����                        ��j�    3      ����3����                        ��j�    4      ����4����                        ��X4_vcswitchX4_vcswitch
 9               `abcSwitches   Generic   X4X4          ������   CParamSubModelType��voltage controlled switch   VCSW{.subckt vcsw 1 2 3 4
S 1 2 3 4 switch
.model switch sw (vt={(Von+Voff)/2} vh={(Von-Voff)/2} ron={Ron} roff={Roff})
.ends   ��  	 CParmDefn    1turnon voltage   ParamSubVon               f�    1turnoff voltage   ParamSubVoffV             f�    0on resistance   ParamSubRonOhm             f�    0off resistance   ParamSubRoffOhm               X #�    ����11      PASA1H�~����#�   ����22      PASA2	   ����#�   ����33      PASA3�8  ����#�   ����44      PASA4�8  ����Switches Generic              8 : `j�   D-      (  D-����                        �� 8  98 	�    �   @      �*   q�   @  `   r 	           	                 D+    	�   D      @  D-��c @            D2     �                   ��                                                           `   D+�                   ��                                                          �   D-�     �       �      ��                                                        �     �   �����     ��                                                        �     �   �����     ��                                                        �     `       �     ��                                                        �    �       �     ��                                                        �     �   �����     ��                                                        �     �       �     ��                                                        � 0   `   �   �    	 ��        	                                               0   `   �   �   0   `   �   �   	[devname]        �������������������������      � 0   �   �   �    
 ��        
                                               0   �   �   �   0   �   �   �   	[refname]       �  �  Y  g  ����   �   <    wxyz{|}    ~          uv �  diode     Miscellaneous      �?       �     � ����        ��������� ���� 27     ��������� ����       ��������� ����       �������� D+D- j�   D+        (  D+����                        ��od1n4007d1n4007    �          �oDiode   Generic   D2D2                D #�    ����D+D+      PASAA��}    #�   ����D-D-      PASAK��}   DiodeDiode	FairchildDO-41             10  j�    M-      ����M-����                        ���	 10 	 510 	�    �    `   `   M+2  	�   s  `   �  M-3   �
  �        IS2    	 �                    ��                                                               M+�                   ��                                                          �   M-�             <     ��                                                        �     �       �     ��                                                        � �����   @   <                  ����                                         ����<   @   �   � ����H   ����t     ��                                                        �  ������� �������  ��          @ @                                           �����x    ��b�����l    
>DA�����l    uT@ @ � ����D   <   |     ��                                                      ����D   <   |   ����D   <   |   [value]       �	  L  �
  �     D   �   |   � ��������B        ��                                                       ��������B      ��������B      	[refname]       f	  b  
       �����      
 ������  ���	   Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       �     � ����    PI��-466.20n      �������� M+M- j�     M+        ����M+����                        ���AmmeterAmmeter   V            ��Analog Meters   Generic   IS2IS2          ����  VAm #�    ����M+M+      PASAM+LVIS����#�   ����M-M-      PASAM-TA
>����Analog MetersAmmeter-verticalGeneric              4  1� j�    L-      ����L-����                        ��� 4  � 4 	�            �   L+K  	�   �   �  �   L-L   @  �          L1     �                    ��                                                           @   L+�                   ��                                                      �   @   L-�� ����,   ���T   
                                                           h   ,   �   T   h   ,   �   T   �   @   h   @           �� ����,  ����T   	                                                           P   ,   h   T   P   ,   h   T   h   @   P   @           �� ����,  ����T                                                              8   ,   P   T   8   ,   P   T   P   @   8   @           �� ����,  ����T                                                                  ,   8   T       ,   8   T   8   @       @           � $   P      X     ��    ���                                                 �    H   $   P     ��                                                        �     P   $   P     ��    ���                                                 �     @       @     ��    (�K	                                                � �   @   �   @     ��       
                                                �     \   �   |     ��                                                           \   �   |       \   �   |   [Inductance]       @  �  �  "      \   �   |   �         �   $     ��                                                               �   $           �   $   	[refname]       @  �  �  +          �   $    ���  �  �  �  ���  �  �  �  �     Inductor     Miscellaneous      �?    
   ��     � ��� {�G�zt?5m      ��������� ���� x     �������� L+L- j�     L+        ����L+����                        ��� Inductor  
 �           ��Passive   Generic   L1L1          ����  L #�    ����L+L+      PASAL+    ����#�   ����L-L-      PASAL-    ����PassiveInductorGeneric              VSource �  j�     1       ����1����                        ��� ��  VSource   s VSource r 	�    {    `       1�  	�   �   �  �   �+   ��   �   	   �                    `   �  2�   `             X1     �                    ��                                                               1�                   ��                                                          �   2�             $     ��    ��)                                                �     \       �     ��                                                        �    8   0   8    	 ��    ��)                                                �     H   @   H     ��    p�Z                                                �     $   @   $     ��                                                       �    \   0   \     ��    D�Z                                                �               ���                                                      �               ���   �Z	                                                � `          $    
 ��        
                                               `          $   `          $   	[devname]        ����������������`          $   � `   $      H     ��                                                       `   $      H   `   $      H   	[refname]       �  �  �  7  `   $      H    ��������    ��    �  �     Battery     Miscellaneous      �?    9 
 Z�     � ����      (@12      �������� 12 �j�    2      ����2����                        ��BatteryBattery
 9 i             ��Sources   Generic   X1X1          ����d���    BATTERY2.SUBCKT Xbattery 1 2
V1 1 2 DC {voltage}
.ENDS
   f�    1battery voltage   ParamSubvoltageV                X #�    ����11      PASA10Ab����#�   ����22      PASA2�1b����SourcesBatteryGeneric              6 p  �j�    M-      ����M-����                        �� 6  o 6 	�    Z    `   �  M+2  	�   �  `   `   M-3   `  �         I_Source    	 �                    ��                                                           �   M+�                   ��                                                              M-�     �       �     ��                                                        �     <             ��                                                        � @   <   �����                  ����                                         ����<   @   �   � ����x   ����L     ��                                                        �  ������� �������  ��          @ @                                           �����H    ��b�����T    
>DA�����T    uT@ @ � ����D   <   |     ��                                                      ����D   <   |   ����D   <   |   [value]       4  l	  ]  �	     D   �   |   � ��������B        ��                                                       ��������B      ��������B      	[refname]       �  �  �  -	     �����      
 ������  ���	   Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       �     � g    @$�$?159.92u      �������� M+M- j�     M+        ����M+����                        ���AmmeterAmmeter   V            ��Analog Meters   Generic   I_SourceI_Source          ����  VAm #�    ����M+M+      PASAM+   @����#�   ����M-M-      PASAM-��W����Analog MetersAmmeter-verticalGeneric              0 >?�    L     �           �   �           �   �               Gnd�	�    �'      @   �.   �       
   �         �                `       Gnd}   �  @          gnd2     �                    ��                                                               Gnd�                   ��     �          AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��     5 (         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��    �׿         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         ����  �     Ground    
Ground DINMiscellaneous      �?       h�       Gnd j�     Gnd        ����Gnd����                        ��gndgnd                 �Analog Meters   Generic   gnd2gnd2          ����  gnd #�    ����GndGnd      GNDAGnd�����SourcesGroundGeneric              0 �   L     0  j�    V-      ����V-����                        ��k ��j�     1       ����1����                        ��j�    4      ����4����                        ��ab  0    J 0 � I m 	�    V        �  1S  	�   �          2T  	�   *   �      3U  	�   R   �   �  4V   �  �         X2     �                    ��                                                           �   1�                   ��                                                          `   2�                   ��                                                      @   `   3�                   ��                                                      @   �   4� @   �   @   �     ��    ��                                                � @   `   @   �     ��                                                        � @   �   @   �    
 ���   ��                                                � H   �   8   �    	 ���   p�H                                                P�    �   �����                  ����                                         �����      �   �����      �   � P   �   0   �               	   ����                                         0   �   P   �   �     `       �     ��       
                                                �    �       �     ��    D�H                                                �     �       �     ��                                                       � 8   �   H   �     ��  � �H        	FIXED_ROT                                        � ,   �      �     ��                                                        � `   �   �   �     ��                                                       `   �   �   �   `   �   �   �   	[refname]       �  �	  2  G
  T   �   �   �   � �   �   @  �     ��                                                       `   `   �   �   `   `   �   �   	[devname]        ����������������T   `   �   �    ������      �  � ��    � �  vcswitch     Miscellaneous      �?   9 
 Z�    � ����      @3      ��������� ����      @3     ��������� ����      �?0.5     ��������� ����    ��.A1meg     �������� 1234 �� j�    3      ����3����                        ���vcswitchvcswitch
 9               �� �Switches   Generic   X2X2          ����d���voltage controlled switch   VCSW{.subckt vcsw 1 2 3 4
S 1 2 3 4 switch
.model switch sw (vt={(Von+Voff)/2} vh={(Von-Voff)/2} ron={Ron} roff={Roff})
.ends   f�    1turnon voltage   ParamSubVon               f�    1turnoff voltage   ParamSubVoffV             f�    0on resistance   ParamSubRonOhm             f�    0off resistance   ParamSubRoffOhm               X #�    ����11      PASA1�S����#�   ����22      PASA2    ����#�   ����33      PASA3�U����#�   ����44      PASA4531E����Switches Generic              VControl @ j�     V+        ����V+����                        ��" 5 G c VControl    VControl �	�    <           V+g  	�   �      �  V-h      �         VCtrl     �                   ��                                                           `   V+�                   ��                                                          �   V-P�     �   �����                   ����                                         �����       �   �����       �   �    �   �����     ��    ��)                                                �     �       �     ��    ��`                                                �     �       �     ��    ��)                                                �     \       �     ��    p�Z                                                � �����   
   �    
 ��               	FIXED_ROT                                        � \   `   \   `     ��                                                      \   `   \   `   \   `   \   `           4  �  4  �                � 0   �   �   �     ��        	                                               0   �   �   �   0   �   �   �   [dc]       �  0	  �  �	          p   @   � 0   \   �   �    	 ��        
                                               0   \   �   �   0   \   �   �   	[refname]       �  �  �  ?	      ����t          !"           �  Voltage Source    Voltage Source DINRoot      �?       ��  CVSourceBehavior     � ����        0      ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       �������� V+V- �volt_sourcevolt_source   +0            �Sources   Generic   VCtrlVCtrl          ����       �0            0      ���������0����      $@10     ���������0            0     ���������0 -1����Mb`?2m     ���������0 -1����Mb`?2m     ���������0�,y�&1�|?7m     ���������0��!
�� �rh�?17m     ��������    �0            0      ���������0����      @5     ���������0����     �f@180     ���������0            0     ���������0            0     ��������    �0            0      ���������0����      �?1     ���������0����      �?1     ���������0            0     ���������0����      �?1     ��������    �0            0      ���������0����      �?1     ���������0            0     ���������0 N  �����>2u     ���������0'  ���ư>1u     ���������0'  ���ư>1u     ��������    �  ���� 0 0      ��������                0      �������� ����       �������� ����       �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������               V #�    ����V+V+      PWR+AV+NDDA����#�   ����V-V-      PWR-AV- � ����Sources Generic              � s N  �o J & 8 � � � =� 5� w 9
 
 
 L  u � � q � ;� 70 # 0                           C � � z � � ) � � � � | ~ � ] [ � W S Q � � � � a Y � _ r�� ; �U < 0 <     �V �             �b      D{ q� � �Z   s� � `  < � B  � � � P � } �� � � y ^ � R X � � * ( : \ � � T � �     ��  CLetter    CEn el model real, els dos inductors estar�n acoplats magn�ticament.  �   }  �      ����Arial����                       Arial     K�   �La tensi� de sortida puja una mica m�s si tenim diodes que converteixen el interruptors en interruptor unidireccionals, que no permeten que la corrent vagi cam a la font.
I la potencia consumida tamb� puja considerablement.�  h  g  i      ����Arial����                       Arial     K�   oLa freq��ncia de traball ha d'estar molt ben ajustada a la freq. de resonancia de les bobines y el condensador.�  5  �  v      ����Arial����                       Arial     K�   ;Ajustant el temps en ON podem ajustar la tensi� de sortida.�  �  J  �      ����Arial����                       Arial     K�   dLa freq��ncia de treball ha de ser lleugerement superior a la corresponent a la freq. de resonancia.�  (  �  i      ����Arial����                       Arial            
 �@ ����        ���������             0     ��������� ����      @5     ���������  ʚ;�������?.1     ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ���� true
     ��������� ����  false     ��������               
                  � ����        ��������� ����       ���������  ����       ���������@ ����       ���������@ ����       ��������               
                  � ����        ��������� ����       ���������@ ����       ���������  ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������               
                 � ����dec     ��������� ����     @�@1k     ��������� ����    ��.A1meg     ��������� ����       20     ��������� ���� true     ��������� ���� true     ��������� ���� true	     ��������� ����  false
     ��������               
                 �  ����        ���������  ����       ���������  ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����  	     ��������� ����  
     ��������               
                  	 � ����        ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������               
                 � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                    �             0      ���������  /hY333333�?150m     ��������� �� �h㈵��>0.01m     ��������� �� �h㈵��>0.01m     ��������� ���� True     ��������� ����  F     ��������� ���� true     ��������� ����  false     ��������               
                 � ����     @�@1K      ���������  ����       ���������  ����       ���������  ����       ��������               
         ��              �  ����        ��������              
                  �  ����        ��������              
                                  
                 �@ ����        ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ���� true	     ��������� ����  false
     ��������� ���� true     ��������� ����  false     ��������               
                 � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                        � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                 � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                 � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                 �@ ����        ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����decade     ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������               
                 � ����        ��������� ����       ���������@ ����       ���������  ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������               
                        � ����dec     ��������� ����     @�@1k     ��������� ����    ��.A1meg     ��������� ����       20     ��������� ����        0     ��������� ����        0     ��������� ���� true	     ��������� ���� true
     ��������� ����      I@50     ��������� ���� true     ��������� ����  false     ��������               
                         / � ���� x'     ���������     �-���q=1E-12     ��������� @B -C��6?1E-4     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x	     ��������� ���� x!     ��������� ����    �  500
     ��������� ���� x     ��������� ����    �  500     ��������� ���� x$     ��������� ���� x$     ��������� ���� x%     ��������� ���� x"     ���������  ���� x*     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x&     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x+     ��������� ���� x,     ��������� ���� x-     ��������� ���� xg     ��������� ���� xf     ��������� ���� xd     ��������� ���� xe     ��������� ���� xh     ��������� ���� xj     ��������� ���� xi     ��������� ���� xk     ��������� ����    e��A1Gl     ���������             0�     ��������� ����      @5�     ��������� ����      @2.5�     ��������� ����      �?.5�     ��������� ����      @4.5�     ��������� 
   ��&�.>1n�     ��������� 
   ��&�.>1n�     ��������� 
   ��&�.>1n�     ��������� 
   ��&�.>1n�     ��������           ��  CPrimitiveModel    d1n4007   �    1�a��%>2.55e-9      ��������� ���� 27     ���������  �/�$��?0.042     ��������� ����      �?1.75     ���������  �  ��v��(�>5.76e-6     ���������     �]}IW�=1.85e-11     ��������� ����      �?0.75     ��������� ����Zd;�O�?0.333     ��������� ���� 1.11	     ��������� ���� 3.0
     ���������      0     ��������� ���� 1     ��������� ���� 0.5     ��������� ����     @�@1000     ��������� � Ǯ���?9.86e-5     ��������     Diode Generic��   CPrimitiveModelType Junction Diode model����DD   f����� 1.0E-14Saturation current    ProcessisAmp0       e     f����� 27!Parameter measurement temperature    ProcesstnomDeg C0     s     f����� 0Ohmic resistance    ProcessrsOhm0      f     f����� 1Emission Coefficient    Processn 0      g     f����� 0Transit Time    Processttsec0     h     f����� 0Junction capacitance    ProcesscjoF0     i     f����� 0     Processcj0F0     i     f����� 1Junction potential    ProcessvjV0      j     f����� 0.5Grading coefficient    Processm 0      k     f����� 1.11Activation energy    ProcessegeV0     	 l     f����� 3.0#Saturation current temperature exp.    Processxti 0     
 m     f����� 0flicker noise coefficient    Processkf 0      t     f����� 1flicker noise exponent    Processaf 0      u     f����� 0.5#Forward bias junction fit parameter    Processfc 0      n     f����� infReverse breakdown voltage    ProcessbvV0      o     f����� 1.0e-3$Current at reverse breakdown voltage    ProcessibvA0      p     f�����  Ohmic conductance    ProcesscondMho     r        D��     �[                Ariald     h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j                   ����            .I                ��  TSignal                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                     i(i_source)       ����                  ��	                     i(is1)       ����                  ��
                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CDCsweep       
 QRSTUVWXYZ               
                       ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                      i(i_source)       ����                  ��	                      i(is1)       ����                  ��
                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACsweep        klmnopqr               
                       ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                     i(i_source)       ����                  ��	                     i(is1)       ����                  ��
                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  �� 
 CTranSweep       ��������               
                       ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                      i(i_source)       ����                  ��	                      i(is1)       ����                  ��
                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACdisto        �����               
                           ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                      i(i_source)       ����                  ��	                      i(is1)       ����                  ��
                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
         �                 ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                      i(i_source)       ����                  ��	                      i(is1)       ����                  ��
                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                          ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                      i(i_source)       ����                  ��	                      i(is1)       ����                  ��
                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                           ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                      i(i_source)       ����                  ��	                      i(is1)       ����                  ��
                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                           ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                      i(i_source)       ����                  ��	                      i(is1)       ����                  ��
                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
         �             	    ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                     i(i_source)       ����                  ��	                     i(is1)       ����                  ��
                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACnoise        stuvwxyz               
                    
    ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                     i(i_source)       ����                  ��	                     i(is1)       ����                  ��
                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  �         �  ����        ���������  ����       ���������  ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����  	     ��������� ����  
     ��������              
                        ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                     i(i_source)       ����                  ��	                     i(is1)       ����                  ��
                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CFourier        ����               
         ��                   ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                     i(i_source)       ����                  ��	                     i(is1)       ����                  ��
                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACpz        	 {|}~����               
                       ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                     i(i_source)       ����                  ��	                     i(is1)       ����                  ��
                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CDCtf         [\]^_               
                       ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                     i(i_source)       ����                  ��	                     i(is1)       ����                  ��
                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CDCsens         `abcdefghij               
                       ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                      i(i_source)       ����                  ��	                      i(is1)       ����                  ��
                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j                  ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                     i(i_source)       ����                  ��	                     i(is1)       ����                  ��
                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CShow         �              
                       ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                     i(i_source)       ����                  ��	                     i(is1)       ����                  ��
                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CShowmod         �              
                       ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                     i(i_source)       ����                  ��	                     i(is1)       ����                  ��
                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  �� 
 CLinearize        �  ����        ��������               
                       ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                     i(i_source)       ����                  ��	                     i(is1)       ����                  ��
                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CParamTranSweep        �������������               
                       ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                     i(i_source)       ����                  ��	                     i(is1)       ����                  ��
                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  �              ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                      i(i_source)       ����                  ��	                      i(is1)       ����                  ��
                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CParamACSweep                        
                       ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                     i(i_source)       ����                  ��	                     i(is1)       ����                  ��
                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CMonteCarlo_op        ����������������������������               
                              ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                     i(i_source)       ����                  ��	                     i(is1)       ����                  ��
                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CMonteCarlo_dc        ����������������������������               
                       ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                      i(i_source)       ����                  ��	                      i(is1)       ����                  ��
                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CMonteCarlo_ac        ����������������������������               
                       ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                     i(i_source)       ����                  ��	                     i(is1)       ����                  ��
                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CMonteCarlo_tran        �������� 	
               
                       ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                      i(i_source)       ����                  ��	                      i(is1)       ����                  ��
                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACsens        !"#$%&'()*+               
                              ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                      i(i_source)       ����                  ��	                      i(is1)       ����                  ��
                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CNetworkAnalysis        ,-./0123456               
                       ����            P               ��                        v(vcontrol)       ����                  ��                       v(3)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                       v(6)       ����                  ��                       v(7)       ����                  ��                       v(8)       ����                  ��                       i(vctrl)       ����                  ��                      i(i_source)       ����                  ��	                      i(is1)       ����                  ��
                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j                  ����            P              33�=           ��   CDigSimResTemplate                ���       ����  ����:�0�yU>20.00n���   ����                       Arial����                       Arial����                       Arial  �   �  �                                ����  ���� ������       ����  ���� ������                 �               ����  �����       200������         0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial      �       �         �     �   �  �  Circuit1                  ����  ��    ��������                                                                                                                                                                                                                                 g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     ��   CPackageAliasSuperPCBStandardDIODE3      �Eagle	DIODE.LBRDO41-7   AC  �Orcad 	DAX2/DO41      �	Ultiboard	L7DIO.l55DIO_DO41              A                  g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �              A    �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            H  �                L C�� �� K TE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                      �  �                �         �  @                  ���                                                  �  @  �     <   �  <     ��                                                        �     |   �  |     ��                                                        �     �   �  �     ��                                                        �     �   �  �     ��                                                        � �      �  4     ��                                                      �      �  4   �      �  4   [title]                                       � �   D   �  t     ��                                                      �   D   �  t   �   D   �  t   [description]                                       � `   �   h  �     ��                                                      `   �   h  �   `   �   h  �   [id]                                       � �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       �      �   8    ��        	                                                   �   8       �   8  Date :       �    8  �                  � �     �  4   	 ��        
                                              �     �  4  �     �  4  [date]                                       �       t   8    
 ��                                                            t   8         t   8   Title :       �      �                  �    L   �   x     ��                                                         L   �   x      L   �   x   Description :       �  �  �   �                  �    �   �   �     ��                                                         �   �   �      �   �   �   ID :       �  �  �  T                  �    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �  L  (                      #$%&'()*+-./01          ,     	title box    Analog Misc      �?    9 
 Z�     �  ����        ���������  ����       ���������  ����       ���������  ����       ���������  ����       ��������        9                                      ����d��� ����     f�            title                f�            description               f�            id               f�            designer               f�            date                           ����            `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                                                                                            2         �  �              � � �                   ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                          �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   
cgs 76         47 80moh5.6 B 1.4988mvrd nmodel MVCTRL.I �     ��                      TIME� # ) time                      ��                        v(3)      v(3)    TIME                 ��                        i(vctrl)� �   i(vctrl)    TIME                 ��                        v(vcontrol)      v(vcontrol)    TIME                 ��    (v(5)-v(9))                   v(Vp)� �   v(Vp)    TIME                 ��                        
v(vsource)      
v(vsource)    TIME                 ��                       i(i_source)�   � i(i_source)    TIME                 ��                       i(is1)  � � i(is1)    TIME                 ��                       i(is2)� �   i(is2)    TIME                 ��    i(i_source)*v(vsource)                   Pin� # )  ����TIME                 ��                        v(9)      v(9)    TIME                           2         �  �           Time  � � �            �
    ����                       Arial����                       Arial                              ����  ����0�̕A�?1.348140e-001����ZP      ����  ��������C�?1.270661e-001��%��K      ����  ������쁆,@1.426271e+001������      ����  ������<�!���-1.607210e+000������                                                                           �                      �                                                                                                                                                                                                                                                                  �  �                                                                                                                                                                                                                                                                              �  �                                                                                                                                                                                                                                                          1m  0                            100   100                                                             1m  0                            100   100                                1m  0                            100   100                                1m  0                            100   100                                                 
                 1m  0                            100   100                            ��   CPartPackage     ��   CPackageg   DO-41�3 pin diode package                                                                                                                                                                                                                                       �         K�     N      ��   CMiniPartPin    ����V+V+     PWR+V+g      P�   ����V-V-     PWR-V-h     voltage_sourcevoltage_source                          P�    ����M+M+     PASM+i      P�   ����M-M-     PASM-j     	voltmeter	voltmeter                          P�    ����11     PAS1�      P�   ����22     PAS2�     BatteryBattery                          P�    ����GndGnd     GNDGnd}      GndGnd                  P�    ����MM       ��������MarkerMarker                  P�    ����GndGnd     GNDGnd}      GndGnd                  P�    ����M+M+     PASM+2      P�   ����M-M-     PASM-3     Ammeter2Ammeter2                          P�    ����11     PAS1S      P�   ����22     PAS2T     P�   ����33     PAS3U     P�   ����44     PAS4V     vcswitchvcswitch                                          P�    ����MM       ��������MarkerMarker                  P�    ����MM       ��������MarkerMarker                  P�    ����L+L+     PASL+K      P�   ����L-L-     PASL-L     InductorInductor                          P�    ����C+C+     PASC+�      P�   ����C-C-     PASC-�     capacitor_genericcapacitor_generic                          P�    ����L+L+     PASL+K      P�   ����L-L-     PASL-L     InductorInductor                          P�    ����11     PAS1S      P�   ����22     PAS2T     P�   ����33     PAS3U     P�   ����44     PAS4V     vcswitchvcswitch                                          P�    ����M+M+     PASM+2      P�   ����M-M-     PASM-3     Ammeter2Ammeter2                          P�    ����M+M+     PASM+2      P�   ����M-M-     PASM-3     Ammeter2Ammeter2                       L P�    ����D+D+     PASA     P�   ����D-D-     PASK      �   ��   CPackagePin 1 D+   AAr� 2 D-   AKDiodeDiode	Fairchild      1n4007 D1n4007D1            diode-21n40071n4007                          P�    ����MM       ��������MarkerMarker               O P�    ����D+D+     PASA     P�   ����D-D-     PASK      9  r� 1 D+   AAr� 2 D-   AKDiodeDiode	Fairchild      1n4007 D1n4007D2            diode-21n40071n4007                                                                                                                                                                                                                                                                                     
m1     8 8 mm l=100u w                        used                             ��    �����Z��� ��                        X�T                                                                                                                                                           `                               �i��    �i��     � ����                        ���                                   �&��0�u .I �   �                         �                                                                                                                                                                                       ���    �����������                            �i��                            ��               �����                        �@�                            �i��    �i�������@
KCTRL                        ���                            ?Q    �?Q�?Q@QXP                        �P                            Ha    �_\PU�_\`\                        c\                            TRL.      
QVI_SOURCE.I                         G5                              �[�    h\��\��\�0]�                        `�X                            ×sA    S1.I Le�7
JL2.I                         G6                              >DAT    .3478332763E-001                        E.I                              
G5    A
G4 =���
G3 5�                        A
>D                            TAB     72492234E-002
MV                         V �    2 2 2 2 d                                                                         