    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz    ��  CPart    �����   �  �  �����   �  �              voltage_source��  CIntPin    ��  CWire    �        �
   /   �   �      /   �   �                  Marker ��  CExtPin    ��  CVertex
      `   ��  CSegment    �6      �                    
        `      M     �  @          Ctrl1     ��   CPin                   ��                                                           `   M��  TLine     P       `     ��    ��                                                ��  TPolygon     ����    ����   ��                                                         ��  TPoint    0        �   @        �    P        �0   @            ��  
 TTextField    �����        ��                                                          �����         �����      	[refname]       �  1  �  �        �   ,               Marker     Miscellaneous      �?    +   ��   CMarkerBehavior     ��  CValue             0.0      �������� M ��  	 TModelPin ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �         �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               " Analog MiscV   Generic   Ctrl1Ctrl1          ����               Ctrl1  v(Ctrl1)  N ��   CPartPin    ����MM       A     ����RootmarkerGeneric              Ctrl1 �        �   /   �   �      /   �   �                  Marker% 	�    �       �   �&   ( �      �   )                       `      MȘ� �  `          Ctrl1     �                   ��                                                           `   M�     P       `     ��                                                        �     ����    ����   ��                                                         �    0        �   @        �    P        �0   @            �    �����        ��                                                          �����         �����      	[refname]       �  Q  �  �        �   ,    -   + 2 ,      Marker     Miscellaneous      �?    +   �     �             0.0      �������� M !� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      3   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               5 Analog MiscV   Generic   Ctrl1Ctrl1          ����               Ctrl1  v(Ctrl1)  N #�    ����MM       A  �����RootmarkerGeneric              Ctrl1 �        �   /   �   �      /   �   �                  Marker7 	�    �      `   �   : �      �   ;                       `      M���� �  @          Ctrl1     �                   ��                                                           `   M�     P       `     ��     �                                                 �     ����    ����   ��                                                         �    0        �   @        �    P        �0   @            �    �����        ��                                                          �����         �����      	[refname]       �  1  �  �        �   ,    ?   = D >      Marker     Miscellaneous      �?    +   �     �             0.0      �������� M !� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      E   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               G Analog MiscV   Generic   Ctrl1Ctrl1          ����               Ctrl1  v(Ctrl1)  N #�    ����MM       A �������RootmarkerGeneric              Ctrl1 �      �       �   �  �      �   �  �              vcswitch�    �     �    L     �           �   �           �   �               GndM 	�    �   �  �   �   �   �  @   Q          P     �   �1   �  �   �   �   �  @   U         T     S      P     �   P �,   `  �   �   �*   `  @   Y          X     W                      `       Gnd}   `  �          gnd1     �                    ��                                                               Gnd�                   ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��    p�Z         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         [ \ ] _   ^      Ground    
Ground DINMiscellaneous      �?       ��   CGroundBehavior       Gnd ��   CBehPin     Gnd        ����Gnd����                        ��gndgnd                 c Analog Meters   Generic   gnd1gnd1          ����  gnd #�    ����GndGnd      GNDAGnd �)����SourcesGroundGeneric              0 K �   L    �           �   �          �   �              Battery�    �    g �    h    �       _   @  �      _   @  �              Ammeter2i �   �    �   l   �       �   �  �      �   �  �              vcswitch�    �    o �   p   �       �   �  �      �   �  �              vcswitch�    L     r 0 q �   �    �    u    �   /   �   �      /   �   �                  Markerv 	�    �&      �   �   y �      �   z                       `      M� �  `          Ctrl2     �                   ��                                                           `   M�     P       `     ��     �                                                 �     ����    ����   ��                                                         �    0        �   @        �    P        �0   @            �    �����        ��                                                          �����         �����      	[refname]       �  Q  �  �        �   ,    ~   | � }      Marker     Miscellaneous      �?    +   �     �             0.0      �������� M !� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     u �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               � Analog MiscV   Generic   Ctrl2Ctrl2          ����               Ctrl2  v(Ctrl2)  N #�    ����MM       A zzzz����RootmarkerGeneric              Ctrl2 �    u    �   /   �   �      /   �   �                  Marker� 	�    �      `   �#   � �!      �   �                       `      Mhz� �  @          Ctrl2     �                   ��                                                           `   M�     P       `     ��                                                        �     ����    ����   ��                                                         �    0        �   @        �    P        �0   @            �    �����        ��                                                          �����         �����      	[refname]       �  1  �  �        �   ,    �   � � �      Marker     Miscellaneous      �?    +   �     �             0.0      �������� M !� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     u �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               � Analog MiscV   Generic   Ctrl2Ctrl2          ����               Ctrl2  v(Ctrl2)  N #�    ����MM       A pH�����RootmarkerGeneric              Ctrl2 �    u    �   /   �   �      /   �   �                  Marker� 	�    �%   @  `   �   � �+   @  �   �                        `      MG5   �  @          Ctrl2     �                   ��                                                           `   M�     P       `     ��    �@
                                                �     ����    ����   ��                                                         �    0        �   @        �    P        �0   @            �    �����        ��                                                          �����         �����      	[refname]       �  1  �  �        �   ,    �   � � �      Marker     Miscellaneous      �?    +   �     �             0.0      �������� M !� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     u �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               � Analog MiscV   Generic   Ctrl2Ctrl2          ����               Ctrl2  v(Ctrl2)  N #�    ����MM       A �����RootmarkerGeneric              Ctrl2 �    u    �   �����   �  �  �����   �  �              voltage_source� �   L    � 0 	�    �           V+g  	�   �'   @  @   �   � �   @  �   �                            �  V-h   @  �         V2     �                   ��                                                           `   V+�                   ��                                                          �   V-��  TEllipse     �   �����                   ����                                         �����       �   �����       �   �    �   �����     ��                                                        �     �       �     ��    1.I                                                 �     �       �     ��    G4                                                  �     \       �     ��    .I                                                 � �����   
   �    
 ��    G3 �        	FIXED_ROT                                        � \   `   \   `     ��                                                      \   `   \   `   \   `   \   `           T  �  T  �                � 0   �   �   �     ��        	                                               0   �   �   �   0   �   �   �   [dc]       �  P    �          p   @   � 0   \   �   �    	 ��        
                                               0   \   �   �   0   \   �   �   	[refname]       �  �  P  T      ����t       �   � � � � � � � �       �     �  �  Voltage Source    Voltage Source DINRoot      �?       ��  CVSourceBehavior     � ����        0      ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       �������� V+V- b�     V+        ����V+����                        ��b�    V-      ����V-����                        ��volt_sourcevolt_source   +0            � � Sources   Generic   V2V2          ����       �0����      @5      ���������0            0     ���������0            0     ���������0��� ����MbP?1m     ���������0��� ����MbP?1m     ���������0���{�G�zt?5m     ���������0 '�~j�t��?12m     ��������    �0            0      ���������0����      @5     ���������0����     ��@10k     ���������0            0     ���������0            0     ��������    �0            0      ���������0����      �?1     ���������0����      �?1     ���������0            0     ���������0����      �?1     ��������    �0            0      ���������0����      �?1     ���������0            0     ���������0 N  �����>2u     ���������0'  ���ư>1u     ���������0'  ���ư>1u     ��������    �  ���� 0 0      ��������                0      �������� ����       �������� ����       �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������               V #�    ����V+V+      PWR+AV+    ����#�   ����V-V-      PWR-AV- �@
����Sources Generic              Ctrl2 t �   u   �       �   �  �      �   �  �              vcswitch�    �    �   �   J 7 � �    �    �       �   �        �   �                Inductor� �   �    �   �   �       �   �  �       �   �  �               R�    p    � 3 � 	�    �   �  �   �$   � �"   `  �   �"   �2   `      �   �   `  `   �         �     � �   �7   @      �        �         �     �!   � �5   `   
    �    �)   `  �              �   �   �   
                       �                    �  �   R+  	�   �      �   �   �3   �
  �   �   �.   �	  �   
       	    �   �0   �
      �
   �   �                      	    �	   	�   �
   
   �   �       
                                           �   R-      �         R     �                    ��                                                       �   @   R+�                   ��                                                          @   R-�    @   $   0     ��    ��)                                                � 0   P   $   0     ��                                                        � 0   P   <   0     ��    ��)                                                � H   P   <   0     ��    p�Z                                                � H   P   T   0     ��                                                       � `   P   h   @     ��    D�Z                                                � �   @   h   @     ��    ��d                                                � `   P   T   0    	 ��    |�f	                                                �    @       @    
 ��    <�b
                                                �     `   �   �     ��                                                           `   �   �       `   �   �   [resistance]           	  �  �	      `   �   �   �         t   $     ��                                                               t   $           t   $   	[refname]          �  H  �          t   $        resistor    resistor DINMiscellaneous      �?       ��  CResistorBehavior     � ����     @@500      ��������� ���� 27     ��������� ����       ��������� ����       �������� R+R- b�     R+        ����R+����                        ��b�    R-      ����R-����                        �� resistor                '(Passive   Generic   RR          ����    R #�    ����R+R+      PASAR+�)����#�   ����R-R-      PASAR-JV1.����Passivedefault resistor, 1KGeneric              6 � �    �    �       �   �  �      �   �  �              	voltmeter+�   p   ,3 	�              M+i  	�   �   �     M-j   �             IV_VRL    
 �                   ��                                                           `   M+�                   ��                                                      �   `   M-�     `       `     ��    ��                                                � �   `   �   `     ��                                                        �    L      \     ��    ��                                                �     T      T     ��    p�H                                                � �   X   �   X     ��               	FIXED_ROT                                        �� 
 TRectangle     <   �   �                   ����                                             <   �   �   � (   D   �   x     ��                                                      (   D   �   x   (   D   �   x   [value]         �  �  b  (   D   �   x   �        �   0    	 ��        	                                                      �   0          �   0   	[refname]          $  `  �         �   0    8  01294  5:6      3
     	voltmeter    voltmeter_smallMiscellaneous      �?       ��   CVoltmeterBehavior     � ����   H	+�-6.29      �������� M+M- b�     M+        ����M+����                        ��b�    M-      ����M-����                        ��	voltmeter	voltmeter   _            >?Analog Meters   Generic   IV_VRLIV_VRL          ����  IVm #�    ����M+M+      PASAM+    ����#�   ����M-M-      PASAM-    ����Analog Meters Generic              6 �    �   �       _   �         _   �                 capacitor_genericB�   p    C3 	�      �  �   C-�  	�          �   C+�      `	          C1     �                   ��                                                       �   @   C-�                   ��                                                          @   C+�     @   @   @      ��    ��                                                � @       @   `     ��                                                        � `       `   `     ��    ��                                                � `   @   �   @     ��    p�H                                                �     `   �   �     ��                                                           `   �   �       `   �   �   [capacitance]          �
  �        `   �   �   �         �   $     ��                                                               �   $           �   $   	[refname]          `	  �   
          �   $    IJKLM    N      GH     	Capacitor     Miscellaneous      �?       ��  CCapacitorBehavior     � '  ����Mbp?4m      ��������� ���� x     ��������� ����       ��������� ����       �������� C+C- b�     C+        ����C+����                        ��b�    C-      ����C-����                        �� 	capacitor    �           UVPassive   Generic   C1C1          ����  C #�    ����C+C+      PASAC+    ����#�   ����C-C-      PASAC-�rR����Passive Generic              6  (>b�    L-      ����L-����                        ��U 6  � 6 	�    �/   �  �   �   �   �  �   �   �   �  �   ^       ]    �   �$   �  `   `        ]    \    [                   �   L+K  	�     �  �   L-L   �  �          L1     �                    ��                                                           @   L+�                   ��                                                      �   @   L-��   TArc h   ,   �   T    
                                                           h   ,   �   T   h   ,   �   T   �   @   h   @           e� P   ,   h   T    	                                                           P   ,   h   T   P   ,   h   T   h   @   P   @           e� 8   ,   P   T                                                               8   ,   P   T   8   ,   P   T   P   @   8   @           e�     ,   8   T                                                                   ,   8   T       ,   8   T   8   @       @           � $   P      X     ��    ��                                                �    H   $   P     ��                                                        �     P   $   P     ��    ��                                                �     @       @     ��    p�H	                                                � �   @   �   @     ��       
                                                �     \   �   |     ��                                                           \   �   |       \   �   |   [Inductance]       �  �  p  �	      \   �   |   �         �   $     ��                                                               �   $           �   $   	[refname]       �  �  P  �          �   $    cdn  m  l  k  jop  i  h  g  f     Inductor     Miscellaneous      �?    
   ��  CInductorBehavior     � ��� ����MbP?1m      ��������� ���� x     �������� L+L- b�     L+        ����L+����                        ��Y Inductor  
  �           uYPassive   Generic   L1L1          ����  L #�    ����L+L+      PASAL+    ����#�   ����L-L-      PASAL-��N����PassiveInductorGeneric              7  b�    2      ����2����                        ��b�     1       ����1����                        ��u 7   � 7 �   l   � 5 � �   L    � 0 	�    a   �   �  1S  	�   �#   �  �   �   �-   �  @   �   �(   �  @   �   ��   �  @   �           �    �    �   ��4   `  @   �   ��   `  �   �           �            ~             �      2T  	�   {          3U  	�   �      `                       �  4V      �        X4     �                    ��                                                       @   �   1�                   ��                                                      @   `   2�                   ��                                                          `   3�                   ��                                                          �   4�     �       �     ��                                                        �     `       �     ��                                                        �     �       �    
 ���                                                       � �����      �    	 ���                                                       �� D   �   <   �                  ����                                         <   �   D   �   <   �   D   �   7�    �   �����               	   ����                                         �����      �   � @   `   @   �     ��        
                                                � 0   �   @   �     ��                                                        � @   �   @   �     ��                                                        �    �   �����     ��  �             	FIXED_ROT                                        �    �   4   �     ��                                                        � `   �   �   �     ��                                                       `   �   �   �   `   �   �   �   	[refname]          |  �        (   t   L   �     �  <    ��                                                       `   `   �   �   `   `   �   �   	[devname]        ����������������       �   (    �������      ��  �������    � �  vcswitch     Miscellaneous      �?   9 
 ��  CParamSubBehavior    � ����������@4.9      ��������� �����������?1.1     ��������� ����      �?0.5     ��������� ����    ��.A1meg     �������� 1234 yb�    2      ����2����                        ��b�    3      ����3����                        ��b�    4      ����4����                        ��X6_vcswitchX6_vcswitch
 9               y���Switches   Generic   X6X6          ������   CParamSubModelType��voltage controlled switch   VCSW{.subckt vcsw 1 2 3 4
S 1 2 3 4 switch
.model switch sw (vt={(Von+Voff)/2} vh={(Von-Voff)/2} ron={Ron} roff={Roff})
.ends   ��  	 CParmDefn    1turnon voltage   ParamSubVon               ��    1turnoff voltage   ParamSubVoffV             ��    0on resistance   ParamSubRonOhm             ��    0off resistance   ParamSubRoffOhm               X #�    ����11      PASA1d   ����#�   ����22      PASA2�2�����#�   ����33      PASA3VA_I����#�   ����44      PASA4G1  ����Switches Generic              Ctrl2  � � �� �  Ctrl2  r Ctrl2 �   L    r 0 	�    Z        �  1S  	�            2T  	�   �   �      3U  	�   �      @                   �   �  4V   `  �         X6     �                    ��                                                           �   1�                   ��                                                          `   2�                   ��                                                      @   `   3�                   ��                                                      @   �   4� @   �   @   �     ��    ��                                                � @   `   @   �     ��                                                        � @   �   @   �    
 ���   ��                                                � H   �   8   �    	 ���   p�H                                                ��    �   �����                  ����                                         �����      �   �����      �   7� P   �   0   �               	   ����                                         0   �   P   �   �     `       �     ��       
                                                �    �       �     ��    D�H                                                �     �       �     ��                                                       � 8   �   H   �     ��  � �H        	FIXED_ROT                                        � ,   �      �     ��                                                        � `   �   �   �     ��                                                       `   �   �   �   `   �   �   �   	[refname]       �  \  �  �      (   t   L   � `   `   �   �     ��                                                       `   `   �   �   `   `   �   �   	[devname]        ����������������       �   (    �������      ��  �������    � �  vcswitch     Miscellaneous      �?   9 
 �  X #�    ����11      PASA1hKS����#�   ����22      PASA2    ����#�   ����33      PASA3    ����#�   ����44      PASA4�XQ����Switches Generic              3 D� - b�     1       ����1����                        ��'?�V 3   n 3 m �      n Ctrl1 �   L    n 0 	�    �        �  1S  	�   �         2T  	�   *   �      3U  	�   �       `                   �   �  4V   `  �         X3     �                    ��                                                           �   1�                   ��                                                          `   2�                   ��                                                      @   `   3�                   ��                                                      @   �   4� @   �   @   �     ��                                                        � @   `   @   �     ��                                                        � @   �   @   �    
 ���                                                       � H   �   8   �    	 ���                                                       ��    �   �����                  ����                                         �����      �   �����      �   7� P   �   0   �               	   ����                                         0   �   P   �   �     `       �     ��    D�H
                                                �    �       �     ��                                                       �     �       �     ��                                                        � 8   �   H   �     ��  �             	FIXED_ROT                                        � ,   �      �     ��                                                        � `   �   �   �     ��                                                       `   �   �   �   `   �   �   �   	[refname]       �  |  �        (   t   L   �     �  <    ��                                                       `   `   �   �   `   `   �   �   	[devname]        ����������������       �   (    �������      ��  �������    � �  vcswitch     Miscellaneous      �?   9 
 ��    � ����������@4.9      ��������� �����������?1.1     ��������� ����      �?0.5     ��������� ����    ��.A1meg     �������� 1234 �xb�    3      ����3����                        ��b�    4      ����4����                        ��vcswitchvcswitch
 9               �x��Switches   Generic   X3X3          ��������voltage controlled switch   VCSW{.subckt vcsw 1 2 3 4
S 1 2 3 4 switch
.model switch sw (vt={(Von+Voff)/2} vh={(Von-Voff)/2} ron={Ron} roff={Roff})
.ends   ��    1turnon voltage   ParamSubVon               ��    1turnoff voltage   ParamSubVoffV             ��    0on resistance   ParamSubRonOhm             ��    0off resistance   ParamSubRoffOhm               X #�    ����11      PASA1    ����#�   ����22      PASA2    ����#�   ����33      PASA3  � ����#�   ����44      PASA4  �����Switches Generic              5 zk  xb�    M-      ����M-����                        ��� 5  j 5 	�    �   �  �   �   ��   �  �   �                       `   �  M+2  	�   �  `   `   M-3   @  �         VA_Ix1    	 �                    ��                                                           �   M+�                   ��                                                              M-�     �       �     ��                                                        �     <             ��                                                        7� @   <   �����                  ����                                         ����<   @   �   � ����x   ����L     ��                                                        �  ������� �������  ��          @ @                                           �����H    ��b�����T    
>DA�����T    uT@ @ � ����D   <   |     ��                                                      ����D   <   |   ����D   <   |   [value]         �    B     D   �   |   � ��������O        ��                                                       ��������O      ��������O      	[refname]       �   �  =  _     �����      
 �����   	   Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       ��   CAmmeterBehavior     � ����   ��")@12.57      �������� M+M- b�     M+        ����M+����                        ���AmmeterAmmeter   V            
�Analog Meters   Generic   VA_Ix1VA_Ix1          ����  VAm #�    ����M+M+      PASAM+8�W����#�   ����M-M-      PASAM-��W����Analog MetersAmmeter-verticalGeneric              4  b�     1       ����1����                        ��
 4   f 4 e 	�    �   `       1�  	�   V   `   �  2�   @  �          X1     �                    ��                                                               1�                   ��                                                          �   2�             $     ��    ��)                                                �     \       �     ��                                                        �    8   0   8    	 ��    ��)                                                �     H   @   H     ��    p�Z                                                �     $   @   $     ��                                                       �    \   0   \     ��    D�Z                                                �               ���                                                      �               ���   �Z	                                                � `          $    
 ��        
                                               `          $   `          $   	[devname]        ����������������`          $   � `   $      H     ��                                                       `   $      H   `   $      H   	[refname]       `  ,  �  �  `   $      H                   Battery     Miscellaneous      �?    9 
 ��     � ����      (@12      �������� 12 b�    2      ����2����                        ��BatteryBattery
 9 i             Sources   Generic   X1X1          ��������    BATTERY2.SUBCKT Xbattery 1 2
V1 1 2 DC {voltage}
.ENDS
   ��    1battery voltage   ParamSubvoltageV                X #�    ����11      PASA10Ab����#�   ����22      PASA2�1b����SourcesBatteryGeneric              0 s �    L     �           �   �           �   �               Gnd#	�    �   `       Gnd}   �  `          gnd2     �                    ��                                                               Gnd�                   ��    ��         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         &'(*  )     Ground    
Ground DINMiscellaneous      �?       `�       Gnd b�     Gnd        ����Gnd����                        ��gndgnd                 ,Analog Meters   Generic   gnd2gnd2          ����  gnd #�    ����GndGnd      GNDAGnd    ����SourcesGroundGeneric              0 ��    L     �	           �   �           �   �               Gnd.	�    �      @            	        `       Gnd}   �  @          gnd3     �                    ��                                                               Gnd�                   ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         2346  5     Ground    
Ground DINMiscellaneous      �?       `�       Gnd b�     Gnd        ����Gnd����                        ��gndgnd                 8Analog Meters   Generic   gnd3gnd3          ����  gnd #�    ����GndGnd      GNDAGnd    ����SourcesGroundGeneric              0 �   L    J 0 �    L     �           �   �           �   �               Gnd;	�    �      �   �%   �      @   ?         >                `       Gnd}   �  �          gnd4     �                    ��                                                               Gnd�                   ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��    D�H         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��    x�W         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��    X��         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         ABCE  D     Ground    
Ground DINMiscellaneous      �?       `�       Gnd b�     Gnd        ����Gnd����                        ��gndgnd                 GAnalog Meters   Generic   gnd4gnd4          ����  gnd #�    ����GndGnd      GNDAGnd    ����SourcesGroundGeneric              0 �   L     0 �    L     �           �   �           �   �               GndJ	�    �   `       Gnd}   �  `          gnd5     �                    ��                                                               Gnd�                   ��    p�H         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��    D�H         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         MNOQ  P     Ground    
Ground DINMiscellaneous      �?       `�       Gnd b�     Gnd        ����Gnd����                        ��gndgnd                 SAnalog Meters   Generic   gnd5gnd5          ����  gnd #�    ����GndGnd      GNDAGnd�����SourcesGroundGeneric              0 {�    L     �           �   �           �   �               GndU	�    �   `       Gnd}   �  @          gnd6     �                    ��                                                               Gnd�                   ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��       0         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��       �         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         XYZ\  [     Ground    
Ground DINMiscellaneous      �?       `�       Gnd b�     Gnd        ����Gnd����                        ��gndgnd                 ^Analog Meters   Generic   gnd6gnd6          ����  gnd #�    ����GndGnd      GNDAGnd��������SourcesGroundGeneric              0 ��    L     �           �   �           �   �               Gnd`	�    �    `       Gnd}   �  �          gnd7     �                    ��                                                               Gnd�                   ��    �@
         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��    KCTR         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         cdeg  f     Ground    
Ground DINMiscellaneous      �?       `�       Gnd b�     Gnd        ����Gnd����                        ��gndgnd                 iAnalog Meters   Generic   gnd7gnd7          ����  gnd #�    ����GndGnd      GNDAGnd    ����SourcesGroundGeneric              0 �  b�    V-      ����V-����                        ���c �,8G� S�^yi  0    J 0 � I :	�    R    �   �  1S  	�   _  �      2T  	�   <          3U  	�   1      �  4V      �        X2     �                    ��                                                       @   �   1�                   ��                                                      @   `   2�                   ��                                                          `   3�                   ��                                                          �   4�     �       �     ��    ��                                                �     `       �     ��                                                        �     �       �    
 ���   ��                                                � �����      �    	 ���   p�H                                                �� D   �   <   �                  ����                                         <   �   D   �   <   �   D   �   7�    �   �����               	   ����                                         �����      �   � @   `   @   �     ��       
                                                � 0   �   @   �     ��    D�H                                                � @   �   @   �     ��                                                       �    �   �����     ��  � �H        	FIXED_ROT                                        �    �   4   �     ��                                                        � T   �   �   �     ��                                                       T   �   �   �   T   �   �   �   	[refname]       �  \  l  �      (   t   L   �     �  <    ��                                                       T   `   �   �   T   `   �   �   	[devname]        ����������������       �   (    pqrsyz|      u}  ~w�{tv    x �  vcswitch     Miscellaneous      �?   9 
 �  X #�    ����11      PASA18 � ����#�   ����22      PASA2�����#�   ����33      PASA3    ����#�   ����44      PASA4�A�����Switches Generic              Ctrl1 �  b�     V+        ����V+����                        ���" 5 G  Ctrl1    Ctrl1 I	�               V+g  	�   @      �  V-h      �         V1     �                   ��                                                           `   V+�                   ��                                                          �   V-��     �   �����                   ����                                         �����       �   �����       �   �    �   �����     ��    ��)                                                �     �       �     ��    ��`                                                �     �       �     ��    ��)                                                �     \       �     ��    p�Z                                                � �����   
   �    
 ��               	FIXED_ROT                                        � \   `   \   `     ��                                                      \   `   \   `   \   `   \   `             �    �                � 0   �   �   �     ��        	                                               0   �   �   �   0   �   �   �   [dc]       �  P  �  �          p   @   � 0   \   �   �    	 ��        
                                               0   \   �   �   0   \   �   �   	[refname]       �  �    T      ����t       �  ��������      �    � �  Voltage Source    Voltage Source DINRoot      �?       ��     � ����        0      ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       �������� V+V- �kvolt_sourcevolt_source   +0            �kSources   Generic   V1V1          ����       �0            0      ���������0����      @5     ���������0            0     ���������0��� ����MbP?1m     ���������0��� ����MbP?1m     ���������0���{�G�zt?5m     ���������0 '�~j�t��?12m     ��������    �0            0      ���������0����      @5     ���������0����     ��@10k     ���������0            0     ���������0            0     ��������    �0            0      ���������0����      �?1     ���������0����      �?1     ���������0            0     ���������0����      �?1     ��������    �0            0      ���������0����      �?1     ���������0            0     ���������0 N  �����>2u     ���������0'  ���ư>1u     ���������0'  ���ư>1u     ��������    �  ���� 0 0      ��������                0      �������� ����       �������� ����       �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������               V #�    ����V+V+      PWR+AV+NDDA����#�   ����V-V-      PWR-AV- � ����Sources Generic              n f � N ,j J $/ <& 8 � w K� V� r � a� C   L  u p l h � � ' # '     �    \^; �W �`Y S 
� � Q � z U ���   � � � ?) 8 5 8 �V >R _* � �P    �: �  � �@  ]�< � � 1�{ ( � � ~a� y � �Z � X �[T � 	� �    ��  CLetter    OLC formen un filtro per obtenir tensi� senoidal a la RL.
fr=1/(2*pi*sqrt(L*C))�  '
        �?����Arial����                       Arial            
 �@ ����        ���������             0     ��������� ����      @5     ���������  ʚ;�������?.1     ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ���� true
     ��������� ����  false     ��������               
                  � ����        ��������� ����       ���������  ����       ���������@ ����       ���������@ ����       ��������               
                  � ����        ��������� ����       ���������@ ����       ���������  ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������               
                 � ����dec     ��������� ����     @�@1k     ��������� ����    ��.A1meg     ��������� ����       20     ��������� ���� true     ��������� ���� true     ��������� ���� true	     ��������� ����  false
     ��������               
                 �  ����        ���������  ����       ���������  ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����  	     ��������� ����  
     ��������               
                  	 � ����        ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������               
                 � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                    �             0      ���������  �/{�G�z�?80m     ��������� @B -C��6?0.1m     ��������� @B -C��6?0.1m     ��������� ���� True     ��������� ����  F     ��������� ���� true     ��������� ����  false     ��������               
                 � ����     @�@1K      ���������  ����       ���������  ����       ���������  ����       ��������               
         ��              �  ����        ��������              
                  �  ����        ��������              
                                  
                 �@ ����        ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ���� true	     ��������� ����  false
     ��������� ���� true     ��������� ����  false     ��������               
                 � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                        � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                 � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                 � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                 �@ ����        ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����decade     ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������               
                 � ����        ��������� ����       ���������@ ����       ���������  ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������               
                        � ����dec     ��������� ����     @�@1k     ��������� ����    ��.A1meg     ��������� ����       20     ��������� ����        0     ��������� ����        0     ��������� ���� true	     ��������� ���� true
     ��������� ����      I@50     ��������� ���� true     ��������� ����  false     ��������               
                         / � ���� x'     ���������     �-���q=1E-12     ��������� @B -C��6?1E-4     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x	     ��������� ���� x!     ��������� ����    �  500
     ��������� ���� x     ��������� ����    �  500     ��������� ���� x$     ��������� ���� x$     ��������� ���� x%     ��������� ���� x"     ���������  ���� x*     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x&     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x+     ��������� ���� x,     ��������� ���� x-     ��������� ���� xg     ��������� ���� xf     ��������� ���� xd     ��������� ���� xe     ��������� ���� xh     ��������� ���� xj     ��������� ���� xi     ��������� ���� xk     ��������� ����    e��A1Gl     ���������             0�     ��������� ����      @5�     ��������� ����      @2.5�     ��������� ����      �?.5�     ��������� ����      @4.5�     ��������� 
   ��&�.>1n�     ��������� 
   ��&�.>1n�     ��������� 
   ��&�.>1n�     ��������� 
   ��&�.>1n�     ��������                 ��                Ariald         � �|p�|����m�|+j      � �|p�|����m�|+j  ��  COpAnal                         
                        ����            2500              
 ��  TSignal                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                      	v(iv_vrl)       ����                  Ӄ                     	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CDCsweep       
 ����������               
                       ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                       	v(iv_vrl)       ����                  Ӄ                      	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CACsweep        ��������               
                       ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                      	v(iv_vrl)       ����                  Ӄ                     	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  �� 
 CTranSweep       ��������               
                       ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                       	v(iv_vrl)       ����                  Ӄ                      	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CACdisto        �����               
                           ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                       	v(iv_vrl)       ����                  Ӄ                      	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  �        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                           ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                       	v(iv_vrl)       ����                  Ӄ                      	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  �        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                           ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                       	v(iv_vrl)       ����                  Ӄ                      	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  �        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                           ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                       	v(iv_vrl)       ����                  Ӄ                      	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  �        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                           ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                       	v(iv_vrl)       ����                  Ӄ                      	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  �        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                       	    ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                      	v(iv_vrl)       ����                  Ӄ                     	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CACnoise        ��������               
                    
    ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                      	v(iv_vrl)       ����                  Ӄ                     	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ^�         �  ����        ���������  ����       ���������  ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����  	     ��������� ����  
     ��������              
                        ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                      	v(iv_vrl)       ����                  Ӄ                     	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CFourier        ����               
         ��                   ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                      	v(iv_vrl)       ����                  Ӄ                     	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CACpz        	 ���������               
                       ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                      	v(iv_vrl)       ����                  Ӄ                     	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CDCtf         �����               
                       ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                      	v(iv_vrl)       ����                  Ӄ                     	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CDCsens         �����������               
                       ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                       	v(iv_vrl)       ����                  Ӄ                      	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j                  ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                      	v(iv_vrl)       ����                  Ӄ                     	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CShow                        
                       ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                      	v(iv_vrl)       ����                  Ӄ                     	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CShowmod                       
                       ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                      	v(iv_vrl)       ����                  Ӄ                     	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  �� 
 CLinearize        �  ����        ��������               
                       ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                      	v(iv_vrl)       ����                  Ӄ                     	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CParamTranSweep        	
               
                       ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                      	v(iv_vrl)       ����                  Ӄ                     	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  �              ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                       	v(iv_vrl)       ����                  Ӄ                      	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CParamACSweep        ������������               
                       ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                      	v(iv_vrl)       ����                  Ӄ                     	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CMonteCarlo_op         !"#$%&'()*               
                              ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                      	v(iv_vrl)       ����                  Ӄ                     	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CMonteCarlo_dc        +,-./0123456789:;<=>?@ABCDEF               
                       ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                       	v(iv_vrl)       ����                  Ӄ                      	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CMonteCarlo_ac        GHIJKLMNOPQRSTUVWXYZ[\]^_`ab               
                       ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                      	v(iv_vrl)       ����                  Ӄ                     	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CMonteCarlo_tran        cdefghijklmnopqrstuvwxyz{|}~               
                       ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                       	v(iv_vrl)       ����                  Ӄ                      	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CACsens        �����������               
                              ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                       	v(iv_vrl)       ����                  Ӄ                      	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CNetworkAnalysis        �����������               
                       ����            P              
 Ӄ                        v(ctrl1)       ����                  Ӄ                       v(ctrl2)       ����                  Ӄ                       v(3)       ����                  Ӄ                       v(5)       ����                  Ӄ                       v(4)       ����                  Ӄ                       v(6)       ����                  Ӄ                       i(v1)       ����                  Ӄ                       	v(iv_vrl)       ����                  Ӄ                      	i(va_ix1)       ����                  Ӄ	                       i(v2)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j                  ����            P                 >           ��   CDigSimResTemplate                ���       ����  ����:�0�yU>20.00n���   ����                       Arial����                       Arial����                       Arial  �   �  �                                ����  ���� ������       ����  ���� ������                 �               ����  �����       200������         0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial      �       �         �     �   �  �  Circuit1                  ����  ��    ��������                                                                                                                                                                                                                                                                                                                                                     �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J P��                H 4� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                      �  �                7�         �  @                  ���                                                  �  @  �     <   �  <     ��                                                        �     |   �  |     ��                                                        �     �   �  �     ��                                                        �     �   �  �     ��                                                        � �      �  4     ��                                                      �      �  4   �      �  4   [title]                                       � �   D   �  t     ��                                                      �   D   �  t   �   D   �  t   [description]                                       � `   �   h  �     ��                                                      `   �   h  �   `   �   h  �   [id]                                       � �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       �      �   8    ��        	                                                   �   8       �   8  Date :       �    H  �                  � �     �  4   	 ��        
                                              �     �  4  �     �  4  [date]                                       �       t   8    
 ��                                                            t   8         t   8   Title :       �       �                  �    L   �   x     ��                                                         L   �   x      L   �   x   Description :       �  �  �  �                  �    �   �   �     ��                                                         �   �   �      �   �   �   ID :       �  �  �  P                  �    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �  \  8                     JKLMNOPQRTUVWX          S     	title box    Analog Misc      �?    9 
 ��     �  ����        ���������  ����       ���������  ����       ���������  ����       ���������  ����       ��������        9                                      �������� ����     ��            title                ��            description               ��            id               ��            designer               ��            date                           ����            `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                                                                                            2         �  �              � � �                   ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                          �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   
cgs 76         47 80moh5.6 ���� � mvrd nmodel             Ӄ                      TIME� # ) time                      Ӄ                        i(v1)� < � i(v1)    TIME                 Ӄ                        v(3)      v(3)    TIME                 Ӄ                      	i(va_ix1)�   � 	i(va_ix1)    TIME                 Ӄ                        v(ctrl1)      v(ctrl1)    TIME                 Ӄ                        v(6)      v(6)    TIME                 Ӄ                        v(ctrl2)      v(ctrl2)    TIME                 Ӄ    (v(6)-v(3))                  	v(IV_VRL)� �   	v(IV_VRL)    TIME                           2         �  �           Time  � � �                   ����                       Arial����                       Arial                              ����  �����z�`?2.035181e-003��G�6      ����  �����z�`?2.035181e-003��G�6      ����  ����1��{��%�-1.075922e+001������      ����  ����1��{��%�-1.075922e+001������                                                                         �                      �                                                      �  �                                                                                                                                                                                                                                                                                                      �  �                                                                                                                                                                      �                      �                                                                                              �  �                                                                                                              �  �                                                                                                                                                                                          1m  0                            100   100                                                             1m  0                            100   100                                1m  0                            100   100                                1m  0                            100   100                                                 
                 1m  0                            100   100                                ��   CMiniPartPin    ����V+V+     PWR+V+g      o�   ����V-V-     PWR-V-h     voltage_sourcevoltage_source                          o�    ����11     PAS1S      o�   ����22     PAS2T     o�   ����33     PAS3U     o�   ����44     PAS4V     vcswitchvcswitch                                          o�    ����11     PAS1�      o�   ����22     PAS2�     BatteryBattery                          o�    ����R+R+     PASR+      o�   ����R-R-     PASR-     RR                          o�    ����GndGnd     GNDGnd}      GndGnd                  o�    ����M+M+     PASM+i      o�   ����M-M-     PASM-j     	voltmeter	voltmeter                          o�    ����M+M+     PASM+2      o�   ����M-M-     PASM-3     Ammeter2Ammeter2                          o�    ����11     PAS1S      o�   ����22     PAS2T     o�   ����33     PAS3U     o�   ����44     PAS4V     vcswitchvcswitch                                          o�    ����GndGnd     GNDGnd}      GndGnd                  o�    ����GndGnd     GNDGnd}      GndGnd                  o�    ����MM       ��������MarkerMarker                  o�    ����GndGnd     GNDGnd}      GndGnd                  o�    ����MM       ��������MarkerMarker                  o�    ����MM       ��������MarkerMarker                  o�    ����V+V+     PWR+V+g      o�   ����V-V-     PWR-V-h     voltage_sourcevoltage_source                          o�    ����MM       ��������MarkerMarker                  o�    ����GndGnd     GNDGnd}      GndGnd                  o�    ����11     PAS1S      o�   ����22     PAS2T     o�   ����33     PAS3U     o�   ����44     PAS4V     vcswitchvcswitch                                          o�    ����GndGnd     GNDGnd}      GndGnd                  o�    ����MM       ��������MarkerMarker                  o�    ����11     PAS1S      o�   ����22     PAS2T     o�   ����33     PAS3U     o�   ����44     PAS4V     vcswitchvcswitch                                          o�    ����MM       ��������MarkerMarker                  o�    ����GndGnd     GNDGnd}      GndGnd                  o�    ����L+L+     PASL+K      o�   ����L-L-     PASL-L     InductorInductor                          o�    ����C+C+     PASC+�      o�   ����C-C-     PASC-�     capacitor_genericcapacitor_generic                                                                                                                                                                       
m1     8 8 mm l=100u w                        used                            �2�    �Q�R�XR��R�                        T�                                                                                                            (f    x=f � �'f                           �(f                            ,�e    �f � ��e                           ��e                                     �  � ���� �                         .I                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       h�    ���������                        ��                            1200    E-002
JV1.I                             G4                                                                                                                                                                                              �$�    h&��&��&� '�                        H)�                            MJ         W X Y [   Z                          DIN                            sist      resistor DIN                                                                                                                                       1200    E-002
JV1.I                             G4                              3 ��    CTRL1     
>ENDD                        -002                             �N    xW�WX�p 4M                        ЮW                                                                                    2 2 2 2 d                                                                                           