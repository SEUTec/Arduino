    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz      ��  CPart       _   �         _   �                 capacitor_generic��  CIntPin    ��  CWire     �      �   ����  �  �  ����  �  �              switch_time�    �    	 �   
   �       _   @  �      _   @  �              Ammeter2�    �    �      �       _   @  �      _   @  �              Ammeter2�    �    �        �           �   �          �   �              Battery �   �     �         �           �   �           �   �               Gnd ��  CExtPin    ��  CVertex+   `  `   ��  CSegment<   �   `  `	                 �+   �J      `   �,   �      �   "         !                 �1    �'   �  `   �   �O   �  `   �    ' �C   @  `   ( �	   ) �   @  `   * �)   �!   @  `   ,          +              �   �<   @  �   .         )              & �/   �L   �  `   0          '          %     $ �   �1   �  �   2         %                          `       Gnd}      `          gnd1     ��   CPin                    ��                                                               Gnd��  TLine                   ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        6�         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        6�    ,   4   ,     ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        6�    8   (   8     ��    p�Z         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         5 7 8 :   9      Ground    
Ground DINMiscellaneous      �?       ��   CGroundBehavior       Gnd ��   CBehPin     Gnd        ����Gnd����                        ��gndgnd                 > Analog Meters   Generic   gnd1gnd1          ����  gnd ��   CPartPin    ����GndGnd      GNDAGnd �)����SourcesGroundGeneric              0  �       �       _   �  �      _   �  �              
Voltmeter2�        B 8 A �    �(          �2   �H      �   F �5   G �A   `  �   �-   I �   `  �   J            H �4   I �M   �  �   �#   M �:   �  @   N             L �&   M �9   �  �   �%   �$   @  �   �   �E   @  �   T �   U �?   @  �   V                S     R �!   S �2   @      X                 Q     P �   Q �)   �  �   Z                                        E                `   `   M+k  �   #   `   �  M-l   �   �          IV_Vx1    
 4�                    ��                                                               M+4�                   ��                                                          �   M-6�     �       �     ��    ��                                                6�             <     ��    
NVA                                                6�    $      4     ��    ��                                                6�    ,      ,     ��    p�H                                                6�    �      �     ��               	FIXED_ROT                                        �� 
 TRectangle     <   �   �                  ����                                             <   �   �   ��  
 TTextField    D   �   x     ��                                                         D   �   x      D   �   x   [value]       �   l  �  �     D   �   x   f� 8      �   0    	 ��        	                                               8      �   0   8      �   0   	[refname]       h  �  �  o  8      �   0    ] ^ a b c e g     h       `   _ 
     Voltemeter-Vert    Voltemeter-Vert_smallMiscellaneous      �?       ��   CVoltmeterBehavior     ��  CValue ����      (@12.00      �������� M+M- =�     M+        ����M+����                        ��=�    M-      ����M-����                        ��	voltmeter	voltmeter   k            m n Analog Meters   Generic   IV_Vx1IV_Vx1          ����  IVm ?�    ����M+M+      PASAM+@������?�   ����M-M-      PASAM-�����Analog MetersVoltmeter-verticalGeneric              0 �         �       �   �         �   �                 1n4007q �   �    �   t     12 �    t    �       �   �         �   �                 1n4007v �      w 8 �    �N   @  �   �3   z �K   @  @   �$   �F   @  @   �.   �@   @  @            ~     } �'   ~ �   @  �	   �6   �   �  �	   �        �     � �   � �I   @  @   �                     �   �"   @  �   �   �-   �  �   �        �     �   �/   @  �   �        �     �     ~         |     { �*   | �    @  @   �                                   @  D+   �   W          D-    @  `         D3     4�                   ��                                                           �   D+4�                   ��                                                          `   D-6� �����       �      ��    ���                                                 6�     �       �     ��                                                        6� �����       �     ��    ���                                                 6�     �       �     ��    (�K                                                6� �����       �     ��                                                       6�     �      �     ��    ��K                                                6�     �       `     ��    ��K                                                f� d   �   $  �    	 ��        	                                               0   `   �   �   0   `   �   �   	[devname]        �������������������������      f� 0   �   �   �    
 ��        
                                               0   �   �   �   0   �   �   �   	[refname]       �    Y  �  ����   �   <    � � � � � � �     � �           � �  �
  diode     Miscellaneous      �?       ��  CDiodeBehavior     k� ����  F      ��������k� ���� x     ��������k� ���� x     ��������k� ���� x     �������� D+D- =�     D+        ����D+����                        ��=�    D-      ����D-����                        ��d1n4007d1n4007    �          � � Diode   Generic   D3D3                D ?�    ����D+D+      PASAA   `����?�   ����D-D-      PASAK��P����DiodeDiode	FairchildDO-41             12 s �   t   �       S   �  ,      S   �  ,              Ammeter�    �    �   �   �       �   �        �   �                Inductor�    �    �    �    �       �   �  �       �   �  �               R� �      � 3 �    �0   @  �	   �;   � �      �	   �                        �  �   R+  �   �   �	  �	   �   �8   �  �	   � �"   �Q   �  @   �:   �G   �  @   � �(   �>   �  �   �        �     �   � �B   �  @   �                 �     �0   � �,   `  @   �            �   �P   �  �   �   � �      �   �             �   �*   �  �   �         �     �     �     �     �     �   � �D   �  @   �                �                  �   R-   �	   	         R     4�                    ��                                                       �   @   R+4�                   ��                                                          @   R-6�    @   $   0     ��    ��)                                                6� 0   P   $   0     ��                                                        6� 0   P   <   0     ��    ��)                                                6� H   P   <   0     ��    p�Z                                                6� H   P   T   0     ��                                                       6� `   P   h   @     ��    D�Z                                                6� �   @   h   @     ��    ��d                                                6� `   P   T   0    	 ��    |�f	                                                6�    @       @    
 ��    <�b
                                                f�     `   �   �     ��                                                           `   �   �       `   �   �   [resistance]       �	   
  `
  �
      `   �   �   f�         t   $     ��                                                               t   $           t   $   	[refname]       �	   	  
  �	          t   $    � � � � � � � � � � � � �    resistor    resistor DINMiscellaneous      �?       ��  CResistorBehavior     k� �������(\��?0.58      ��������k� ���� 27     ��������k� ����       ��������k� ����       �������� R+R- =�     R+        ����R+����                        ��=�    R-      ����R-����                        �� resistor                � � Passive   Generic   RR          ����    R ?�    ����R+R+      PASAR+JV1.����?�   ����R-R-      PASAR-�)����Passivedefault resistor, 1KGeneric              5 �  � =�     L+        ����L+����                        �� 5   � 5 � �    �        �   L+K  �   �   �  �	   �9   � �.   @  �	   �                      �  �   L-L       	          L1     4�                    ��                                                           @   L+4�                   ��                                                      �   @   L-��   TArc h   ,   �   T    
                                                           h   ,   �   T   h   ,   �   T   �   @   h   @           � P   ,   h   T    	                                                           P   ,   h   T   P   ,   h   T   h   @   P   @           � 8   ,   P   T                                                               8   ,   P   T   8   ,   P   T   P   @   8   @           �     ,   8   T                                                                   ,   8   T       ,   8   T   8   @       @           6� $   P      X     ��    ��                                                6�    H   $   P     ��     �                                                  6�     P   $   P     ��    ��                                                6�     @       @     ��    p�H	                                                6� �   @   �   @     ��       
                                                f�     \   �   |     ��                                                           \   �   |       \   �   |   [Inductance]          
  �  �
      \   �   |   f�         �   $     ��                                                               �   $           �   $   	[refname]           	  r  �	          �   $    � � �   �   �   �   � � �   �   �   �   �      Inductor     Miscellaneous      �?    
   ��  CInductorBehavior     k� ��� �������?100m      ��������k� ���� x     �������� L+L- � =�    L-      ����L-����                        �� Inductor  
              � � Passive   Generic   L1L1          ����  L ?�    ����L+L+      PASAL+������?�   ����L-L-      PASAL-P������PassiveInductorGeneric              16 �  � =�     M+        ����M+����                        �� 16   � 16 � �    �        �   M+0  �   �   �  �   M-1   @   	          VA_IL    	 4�                   ��                                                           @   M+4�                   ��                                                      �   @   M-6� �   @   �   @     ��    ��                                                6�     @       @     ��                                                        6� 4   X   `   X     ��    ��                                                d�        �   d                   ����                                                �   d   ��  TPolygon ����������������  ��          @ @                                           ��  TPointd   X    IX1.�X   P        �X   `    0000@ @ f� $   $   �   L     ��                                                      $   $   �   L   $   $   �   L   [value]       �  l	  �  �	  $   $   �   L   f�     �����        ��                                                           �����          �����      	[refname]       �  �  �  �	      �����         �        	     Ammeter    Ammeter_smallMiscellaneous      �?       ��   CAmmeterBehavior     k� ����   `��9�-6.05n      �������� M+M- � =�    M-      ����M-����                        ��AmmeterAmmeter   �            � Analog Meters   Generic   VA_ILVA_IL          ����  VAm ?�    ����M+M+      PASAM+0�M����?�   ����M-M-      PASAM- ������Analog MetersAmmeterGeneric              12 �    t    �   ����  �  �  ����  �  �              switch_time�       0 �    �        �  SW+=  �   /          SW->   @  �	         X2    
 4�                   ��                                                           �   SW+4�                    ��                                                             SW-� �����                                                                      ����|       �   ����|       �       �       �           6�     �       �     ��    ���                                                 6�     �       �     ��    `                                                   6�     �            ��    ���                                                 6� (   �       �     ��    (�K                                                6�     �      �     ��                                                       f� 8   �   �   �     ��                                                       8   �   �   �   8   �   �   �   	[refname]       �  �  Z  {         t   @   f� 8   |   �   �    	 ��        	                                               8   |   �   �   8   |   �   �   	[devname]        ����������������    �����            !  
 �  Switch_Open     Miscellaneous      �?   9 
 ��  CParamSubBehavior    k� @T� ��H�}M?0.9m      ��������k�  ��{�G�z�?10m     ��������k� ����      �?0.5     ��������k� ����    ��.A1meg     �������� 45 =�     4       ����4����                        ��=�    5      ����5����                        ��X2_switch_timeX2_switch_time
 9 V            ()Switches   Generic   X2X2          ������   CParamSubModelType��time controlled switch   TIME_SWITCH�.subckt tswitch 4 5
S 4  5  3 0 switch
V0 3  0 DC 0 PWL ( 0 0
+ {time_on-.000000001} 0
+ {time_on+.000000001}  1
+ {time_off-.000000001} 1
+ {time_off+.000000001} 0)

IVm0 3  0 0

.model switch SW  vt = .5   vh = 0   ron = {res_on}   roff = {res_off}  
.ends   ��  	 CParmDefn     time the switch closes   ParamSubtime_ons              ,�    1time the switch opens   ParamSubtime_offs             ,�    1resistance when switch closed   ParamSubres_onOhm             ,�    1megresistance when switch open   ParamSubres_offOhm               X ?�    ����SW+4      PASASW+������?�   ����SW-5      PASASW-   �����SwitchesTime Controlled SwitchGeneric              12 �   t   �       �   �  �      �   �  �              	voltmeter�        43 3�    �           M+i  �   �   �     M-j      �          IV_VL    
 4�                   ��                                                           `   M+4�                   ��                                                      �   `   M-6�     `       `     ��    ��                                                6� �   `   �   `     ��                                                        6�    L      \     ��    ��                                                6�     T      T     ��    p�H                                                6� �   X   �   X     ��               	FIXED_ROT                                        d�     <   �   �                   ����                                             <   �   �   f� (   D   �   x     ��                                                      (   D   �   x   (   D   �   x   [value]       x  l  �  �  (   D   �   x   f�        �   0    	 ��        	                                                      �   0          �   0   	[refname]       `  �  ~  o         �   0    ?  89:@<  =A>      ;
     	voltmeter    voltmeter_smallMiscellaneous      �?       i�     k� *}��      ��-29.56u      �������� M+M- =�     M+        ����M+����                        ��=�    M-      ����M-����                        ��	voltmeter	voltmeter   _            DEAnalog Meters   Generic   IV_VLIV_VL          ����  IVm ?�    ����M+M+      PASAM+    ����?�   ����M-M-      PASAM-    ����Analog Meters Generic              12 �   t   �   ����  �  �  ����  �  �              switch_time�        I8 H�    Y        �  SW+=  �   �          SW->   @  �         X3    
 4�                   ��                                                           �   SW+4�                    ��                                                             SW-� �����                                                                      ����|       �   ����|       �       �       �           6�     �       �     ��    ���                                                 6�     �       �     ��                                                        6�     �            ��    ���                                                 6� (   �       �     ��    (�K                                                6�     �      �     ��                                                       f� 8   �   �   �     ��                                                       8   �   �   �   8   �   �   �   	[refname]       �  �  Z  [         t   @   f� 8   |   �   �    	 ��        	                                               8   |   �   �   8   |   �   �   	[devname]        ����������������    �����       N  PQRMT  UVS  O
 �  Switch_Open     Miscellaneous      �?   9 
 "�    k�  h�	����Mb�?16m      ��������k�  ��{�G�z�?20m     ��������k� ����      �?0.5     ��������k� ����    ��.A1meg     �������� 45 =�     4       ����4����                        ��=�    5      ����5����                        ��X4_switch_timeX4_switch_time
 9 ^�            \]Switches   Generic   X3X3          ����*���time controlled switch   TIME_SWITCH�.subckt tswitch 4 5
S 4  5  3 0 switch
V0 3  0 DC 0 PWL ( 0 0
+ {time_on-.000000001} 0
+ {time_on+.000000001}  1
+ {time_off-.000000001} 1
+ {time_off+.000000001} 0)

IVm0 3  0 0

.model switch SW  vt = .5   vh = 0   ron = {res_on}   roff = {res_off}  
.ends   ,�     time the switch closes   ParamSubtime_ons              ,�    1time the switch opens   ParamSubtime_offs             ,�    1resistance when switch closed   ParamSubres_onOhm             ,�    1megresistance when switch open   ParamSubres_offOhm               X ?�    ����SW+4      PASASW+X2.I����?�   ����SW-5      PASASW- @A
����SwitchesTime Controlled SwitchGeneric              12  =�    C-      ����C-����                        ��E=�    D-      ����D-����                        ��]� ( 12  r 12 �    -        @  D+   �   �          D-    @   
         D2     4�                   ��                                                           �   D+4�                   ��                                                          `   D-6� �����       �      ��    ���                                                 6�     �       �     ��                                                        6� �����       �     ��    ���                                                 6�     �       �     ��    (�K                                                6� �����       �     ��                                                       6�     �      �     ��    ��K                                                6�     �       `     ��    ��K                                                f� d   �   $  �    	 ��        	                                               0   `   �   �   0   `   �   �   	[devname]        �������������������������      f� 0   �   �   �    
 ��        
                                               0   �   �   �   0   �   �   �   	[refname]       �  �  Y  �  ����   �   <    klmnopq    rs          ij �
  diode     Miscellaneous      �?       ��     k� ����  F      ��������k� ���� x     ��������k� ���� x     ��������k� ���� x     �������� D+D- =�     D+        ����D+����                        ��fd1n4007d1n4007               yfDiode   Generic   D2D2                D ?�    ����D+D+      PASAA�
MV����?�   ����D-D-      PASAK 
G9����DiodeDiode	FairchildDO-41             0 �         �       �   �         �   �                 1n4007|�      }3 �    1        @  D+   �   �          D-    �   
         D4     4�                   ��                                                           �   D+4�                   ��                                                          `   D-6� �����       �      ��    ���                                                 6�     �       �     ��                                                        6� �����       �     ��    ���                                                 6�     �       �     ��                                                       6� �����       �     ��    ��K                                                6�     �      �     ��    ��K                                                6�     �       `     ��                                                        f� d   �   $  �    	 ��        	                                               0   `   �   �   0   `   �   �   	[devname]        �������������������������      f� 0   �   �   �    
 ��        
                                               0   �   �   �   0   �   �   �   	[refname]       0	  �  �	  �  ����   �   <    �������    ��          �� �
  diode     Miscellaneous      �?       ��     k� ����  F      ��������k� ���� x     ��������k� ���� x     ��������k� ���� x     �������� D+D- =�     D+        ����D+����                        ��=�    D-      ����D-����                        ��d1n4007d1n4007    @          ��Diode   Generic   D4D4                D ?�    ����D+D+      PASAA    ����?�   ����D-D-      PASAK    ����DiodeDiode	FairchildDO-41             0 �       �   ����  �  �  ����  �  �              switch_time�        �3 ��    �        �  SW+=  �   3          SW->   �  �	         X4    
 4�                   ��                                                           �   SW+4�                    ��                                                             SW-� �����                                                                      ����|       �   ����|       �       �       �           6�     �       �     ��    ���                                                 6�     �       �     ��                                                        6�     �            ��    ���                                                 6� (   �       �     ��    (�K                                                6�     �      �     ��                                                       f� 8   �   �   �     ��                                                       8   �   �   �   8   �   �   �   	[refname]       H  �  �  {         t   @   f� 8   |   �   �    	 ��        	                                               8   |   �   �   8   |   �   �   	[devname]        ����������������    �����       �  �����  ���  �
 �  Switch_Open     Miscellaneous      �?   9 
 "�    k�  h�	����Mb�?16m      ��������k� ����������?25m     ��������k� ����      �?0.5     ��������k� ����    ��.A1meg     �������� 45 =�     4       ����4����                        ��=�    5      ����5����                        ��X3_switch_time_0X3_switch_time_0
 9  @            ��Switches   Generic   X4X4          ����*���time controlled switch   TIME_SWITCH�.subckt tswitch 4 5
S 4  5  3 0 switch
V0 3  0 DC 0 PWL ( 0 0
+ {time_on-.000000001} 0
+ {time_on+.000000001}  1
+ {time_off-.000000001} 1
+ {time_off+.000000001} 0)

IVm0 3  0 0

.model switch SW  vt = .5   vh = 0   ron = {res_on}   roff = {res_off}  
.ends   ,�     time the switch closes   ParamSubtime_ons              ,�    1time the switch opens   ParamSubtime_offs             ,�    1resistance when switch closed   ParamSubres_onOhm             ,�    1megresistance when switch open   ParamSubres_offOhm               X ?�    ����SW+4      PASASW+�ȶ
����?�   ����SW-5      PASASW-zzzz����SwitchesTime Controlled SwitchGeneric              0  =�    2      ����2����                        ��> y�n �)  0    0 �    �   `  �   �7   �   `  @   �        �               `       1�  �      `   �  2�      �          XBattery     4�                    ��                                                               14�                   ��                                                          �   26�             $     ��    ��)                                                6�     \       �     ��                                                        6�    8   0   8    	 ��    ��)                                                6�     H   @   H     ��    p�Z                                                6�     $   @   $     ��                                                       6�    \   0   \     ��    D�Z                                                6�               ���                                                      6�               ���   �Z	                                                f� `          $    
 ��        
                                               `          $   `          $   	[devname]        ����������������`          $   f� :   �����   ����  ��                                                       :   �����   ����:   �����   ����	[refname]       �  \  I    `   $      H    ��������    ��    �  �     Battery     Miscellaneous      �?    9 
 "�     k� ����      (@12      �������� 12 =�     1       ����1����                        ���BatteryBattery
 9 i             ��Sources   Generic   XBatteryXBattery          ����*���    BATTERY2.SUBCKT Xbattery 1 2
V1 1 2 DC {voltage}
.ENDS
   ,�    1battery voltage   ParamSubvoltageV                X ?�    ����11      PASA1�1b����?�   ����22      PASA20Ab����SourcesBatteryGeneric              4   �=�     M+        ����M+����                        �� 4    4  �    �   `   �  M+2  �   K   `   `   M-3      `         VA_Ix1    	 4�                    ��                                                           �   M+4�                   ��                                                              M-6�     �       �     ��                                                        6�     <             ��                                                        d� @   <   �����                  ����                                         ����<   @   �   6� ����x   ����L     ��                                                        �  ������� �������  ��          @ @                                           �����H    ��b�����T    
>DA�����T    uT@ @ f� ����D   <   |     ��                                                      ����D   <   |   ����D   <   |   [value]       �  ,  �  �     D   �   |   f� ��������O        ��                                                       ��������O      ��������O      	[refname]       �  ?    �     �����      
 ������  ���	   Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       �     k� �Hl9   @���?96.34m      �������� M+M- �=�    M-      ����M-����                        ��AmmeterAmmeter   V            ��Analog Meters   Generic   VA_Ix1VA_Ix1          ����  VAm ?�    ����M+M+      PASAM+��W����?�   ����M-M-      PASAM-8�W����Analog MetersAmmeter-verticalGeneric              8 C  x J�      �       �   �         �   �                 1n4007�        �3 ��    �        @  D+   �   [          D-    �  `         D1     4�                   ��                                                           �   D+4�                   ��                                                          `   D-6� �����       �      ��    ���                                                 6�     �       �     ��                                                        6� �����       �     ��    ���                                                 6�     �       �     ��                                                       6� �����       �     ��    ��K                                                6�     �      �     ��    ��K                                                6�     �       `     ��    10                                                  f� d   �   $  �    	 ��        	                                               0   `   �   �   0   `   �   �   	[devname]        �������������������������      f� 0   �   �   �    
 ��        
                                               0   �   �   �   0   �   �   �   	[refname]       0	    �	  �  ����   �   <    �������    ��          �� �
  diode     Miscellaneous      �?       ��     k� ����  F      ��������k� ���� x     ��������k� ���� x     ��������k� ���� x     �������� D+D- =�     D+        ����D+����                        ��=�    D-      ����D-����                        ��d1n4007d1n4007   ^�          ��Diode   Generic   D1D1                D ?�    ����D+D+      PASAAA
G5����?�   ����D-D-      PASAKG7  ����DiodeDiode	FairchildDO-41             8  ��\m � =�     M+        ����M+����                        �� 8    8  �    O    `   `   M+2  �   �7   �  �   �8   ��#   �      �                     `   �  M-3   @  �          VA_X1    	 4�                    ��                                                               M+4�                   ��                                                          �   M-6�             <     ��    x�R                                                6�     �       �     ��     zT                                                d�     <   �   �                  ����                                             <   �   �   6� �   H   �   t     ��    (�K                                                � ����������������  ��          @ @                                           ��   x    h�P��   l    �  ��   l        @ @ f�    D   �   |     ��                                                         D   �   |      D   �   |   [value]       L  �  1  :     D   �   |   f� D   ����       ��                                                       D   ����     D   ����     	[refname]         �  A  j     �����      
 ��   		     Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       �     k� ,�     �N@�> 6.02u      �������� M+M- �=�    M-      ����M-����                        ��AmmeterAmmeter   �            �Analog Meters   Generic   VA_X1VA_X1          ����  VAm ?�    ����M+M+      PASAM+PǕ����?�   ����M-M-      PASAM-�������Analog MetersAmmeter-verticalGeneric              15  =�     4       ����4����                        �� 15    15  �    �       �  SW+=  �   �          SW->   �  �         X1    
 4�                   ��                                                           �   SW+4�                    ��                                                             SW-� �����                                                                      ����|       �   ����|       �       �       �           6�     �       �     ��    ���                                                 6�     �       �     ��                                                        6�     �            ��    ���                                                 6� (   �       �     ��    (�K                                                6�     �      �     ��                                                       f� 8   �   �   �     ��                                                       8   �   �   �   8   �   �   �   	[refname]       H  �  �  [         t   @   f� 8   |   �   �    	 ��        	                                               8   |   �   �   8   |   �   �   	[devname]        ����������������    �����             
 �  Switch_Open     Miscellaneous      �?   9 
 "�    k� ��� ����MbP?1m      ��������k� ���{�G�zt?5m     ��������k� ����      �?0.5     ��������k� ����    ��.A1meg     �������� 45 =�    5      ����5����                        ��switch_timeswitch_time
 9               !Switches   Generic   X1X1          ����*���time controlled switch   TIME_SWITCH�.subckt tswitch 4 5
S 4  5  3 0 switch
V0 3  0 DC 0 PWL ( 0 0
+ {time_on-.000000001} 0
+ {time_on+.000000001}  1
+ {time_off-.000000001} 1
+ {time_off+.000000001} 0)

IVm0 3  0 0

.model switch SW  vt = .5   vh = 0   ron = {res_on}   roff = {res_off}  
.ends   ,�     time the switch closes   ParamSubtime_ons              ,�    1time the switch opens   ParamSubtime_offs             ,�    1resistance when switch closed   ParamSubres_onOhm             ,�    1megresistance when switch open   ParamSubres_offOhm               X ?�    ����SW+4      PASASW+    ����?�   ����SW-5      PASASW-    ����SwitchesTime Controlled SwitchGeneric              3 �5�� ~ =�     C+        ����C+����                        ��� D��!� 3   3 u �    �   �  �   C-�  �   �        �   C+�   `  �          C1     4�                   ��                                                       �   @   C-4�                   ��                                                          @   C+6�     @   @   @      ��    ���                                                 6� @       @   `     ��    �b�                                                6� `       `   `     ��    ���                                                 6� `   @   �   @     ��    (�K                                                f�     `   �   �     ��                                                           `   �   �       `   �   �   [capacitance]       `  �  �  .	      `   �   �   f�         �   $     ��                                                               �   $           �   $   	[refname]       `  �  �  +          �   $    ./012    3      ,-     	Capacitor     Miscellaneous      �?       ��  CCapacitorBehavior     k� '  �dy���=20p      ��������k� ���� x     ��������k� ����       ��������k� ����       �������� C+C- )e 	capacitor                )ePassive   Generic   C1C1          ����  C ?�    ����C+C+      PASAC+�R����?�   ����C-C-      PASAC-P�����Passive Generic               �  4                   r �I�     � � B w }       t   �  
 � = . =                 � *         2 &   T   Z   � � � V � . � � � � � ( X � N } R P � � , �   " J  0 � $ F { L H � ��� � �  R 6 R                              �   �  � �   �    � # + �   K � � - � �S     % E [ �  � � � � � 3 Y         �� Q O   /   � W � I � ) � U ~ � G � ! | 1 M z ' � �    ��  CLetter    �Los dos interruptores se ponen en ON al mismo tiempo.
X2 se pone en OFF, deja de fluir corriente desde la fuente.
X3 sigue en ON, por donde circula la corriente adem�s de por D2.
X3 passa a OFF, entonces la corriente retorna a la fuente a trav�s de D1 y D2.
�   2  �  S  -����Arial����                       Arial            
 k�@ ����        ��������k�             0     ��������k� ����      @5     ��������k�  ʚ;�������?.1     ��������k�@ ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ���� true
     ��������k� ����  false     ��������               
                  k� ����        ��������k� ����       ��������k�  ����       ��������k�@ ����       ��������k�@ ����       ��������               
                  k� ����        ��������k� ����       ��������k�@ ����       ��������k�  ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������               
                 k� ����dec     ��������k� ����     @�@1k     ��������k� ����    ��.A1meg     ��������k� ����       20     ��������k� ���� true     ��������k� ���� true     ��������k� ���� true	     ��������k� ����  false
     ��������               
                 k�  ����        ��������k�  ����       ��������k�  ����       ��������k� ����dec     ��������k� ����       ��������k� ����       ��������k� ����  	     ��������k� ����  
     ��������               
                  	 k� ����        ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������               
                 k� ����        ��������k� ����       ��������k� ����       ��������k� ����dec     ��������k� ����       ��������               
                    k�             0      ��������k�  �����Q��?30m     ��������k� �� �h㈵��>0.01m     ��������k� �� �h㈵��>0.01m     ��������k� ���� True     ��������k� ����  F     ��������k� ���� true     ��������k� ����  false     ��������               
                 k� ����     @�@1K      ��������k�  ����       ��������k�  ����       ��������k�  ����       ��������               
         ��              k�  ����        ��������              
                  k�  ����        ��������              
                                  
                 k�@ ����        ��������k�@ ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ���� true	     ��������k� ����  false
     ��������k� ���� true     ��������k� ����  false     ��������               
                 k� ����       5      ��������k� ����       5     ��������k� ����       5     ��������k� ����       5     ��������k� ����       ��������k� ����  	     ��������k� ����  
     ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ���� true     ��������k�@ ����       ��������k�@ ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����dec     ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ���� true     ��������k� ���� true     ��������k� ���� true     ��������k� ����  false     ��������k� ���� true     ��������k� ����  false      ��������k� ���� true!     ��������k� ����  false"     ��������               
                        k� ����       5      ��������k� ����       5     ��������k� ����       5     ��������k� ����       5     ��������k� ����       ��������k� ����  	     ��������k� ����  
     ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ���� true     ��������k�@ ����       ��������k�@ ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����dec     ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ���� true     ��������k� ���� true     ��������k� ���� true     ��������k� ����  false     ��������k� ���� true     ��������k� ����  false      ��������k� ���� true!     ��������k� ����  false"     ��������               
                 k� ����       5      ��������k� ����       5     ��������k� ����       5     ��������k� ����       5     ��������k� ����       ��������k� ����  	     ��������k� ����  
     ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ���� true     ��������k�@ ����       ��������k�@ ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����dec     ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ���� true     ��������k� ���� true     ��������k� ���� true     ��������k� ����  false     ��������k� ���� true     ��������k� ����  false      ��������k� ���� true!     ��������k� ����  false"     ��������               
                 k� ����       5      ��������k� ����       5     ��������k� ����       5     ��������k� ����       5     ��������k� ����       ��������k� ����  	     ��������k� ����  
     ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ���� true     ��������k�@ ����       ��������k�@ ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����dec     ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ���� true     ��������k� ���� true     ��������k� ���� true     ��������k� ����  false     ��������k� ���� true     ��������k� ����  false      ��������k� ���� true!     ��������k� ����  false"     ��������               
                 k�@ ����        ��������k�@ ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����decade     ��������k� ���� true     ��������k� ���� true     ��������k� ���� true     ��������k� ����  false     ��������               
                 k� ����        ��������k� ����       ��������k�@ ����       ��������k�  ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������k� ����       ��������               
                        k� ����dec     ��������k� ����     @�@1k     ��������k� ����    ��.A1meg     ��������k� ����       20     ��������k� ����        0     ��������k� ����        0     ��������k� ���� true	     ��������k� ���� true
     ��������k� ����      I@50     ��������k� ���� true     ��������k� ����  false     ��������               
                         / k� ���� x'     ��������k�     �-���q=1E-12     ��������k� @B -C��6?1E-4     ��������k� ���� x     ��������k� ���� x     ��������k� ���� x     ��������k� ���� x     ��������k� ���� x     ��������k� ���� x     ��������k� ���� x	     ��������k� ���� x!     ��������k� ����    �  500
     ��������k� ���� x     ��������k� ����    �  500     ��������k� ���� x$     ��������k� ���� x$     ��������k� ���� x%     ��������k� ���� x"     ��������k�  ���� x*     ��������k� ���� x     ��������k� ���� x     ��������k� ���� x     ��������k� ���� x&     ��������k� ���� x     ��������k� ���� x     ��������k� ���� x     ��������k� ���� x+     ��������k� ���� x,     ��������k� ���� x-     ��������k� ���� xg     ��������k� ���� xf     ��������k� ���� xd     ��������k� ���� xe     ��������k� ���� xh     ��������k� ���� xj     ��������k� ���� xi     ��������k� ���� xk     ��������k� ����    e��A1Gl     ��������k�             0�     ��������k� ����      @5�     ��������k� ����      @2.5�     ��������k� ����      �?.5�     ��������k� ����      @4.5�     ��������k� 
   ��&�.>1n�     ��������k� 
   ��&�.>1n�     ��������k� 
   ��&�.>1n�     ��������k� 
   ��&�.>1n�     ��������           ��  CPrimitiveModel    d1n4007   k�    1�a��%>2.55e-9      ��������k� ���� 27     ��������k�  �/�$��?0.042     ��������k� ����      �?1.75     ��������k�  �  ��v��(�>5.76e-6     ��������k�     �]}IW�=1.85e-11     ��������k� ����      �?0.75     ��������k� ����Zd;�O�?0.333     ��������k� ���� 1.11	     ��������k� ���� 3.0
     ��������k�      0     ��������k� ���� 1     ��������k� ���� 0.5     ��������k� ����     @�@1000     ��������k� � Ǯ���?9.86e-5     ��������     Diode Generic��   CPrimitiveModelType Junction Diode model����DD   ,����� 1.0E-14Saturation current    ProcessisAmp0       e     ,����� 27!Parameter measurement temperature    ProcesstnomDeg C0     s     ,����� 0Ohmic resistance    ProcessrsOhm0      f     ,����� 1Emission Coefficient    Processn 0      g     ,����� 0Transit Time    Processttsec0     h     ,����� 0Junction capacitance    ProcesscjoF0     i     ,����� 0     Processcj0F0     i     ,����� 1Junction potential    ProcessvjV0      j     ,����� 0.5Grading coefficient    Processm 0      k     ,����� 1.11Activation energy    ProcessegeV0     	 l     ,����� 3.0#Saturation current temperature exp.    Processxti 0     
 m     ,����� 0flicker noise coefficient    Processkf 0      t     ,����� 1flicker noise exponent    Processaf 0      u     ,����� 0.5#Forward bias junction fit parameter    Processfc 0      n     ,����� infReverse breakdown voltage    ProcessbvV0      o     ,����� 1.0e-3$Current at reverse breakdown voltage    ProcessibvA0      p     ,�����  Ohmic conductance    ProcesscondMho     r        D��     �#W�                Ariald     ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  COpAnal                         
                        ����                              ��  TSignal                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                      v(iv_vl)       ����                  y�                     	i(va_ix1)       ����                  y�                     i(x4)       ����                  y�                     i(va_il)       ����                  y�                      	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CDCsweep       
 >?@ABCDEFG               
                       ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                       v(iv_vl)       ����                  y�                      	i(va_ix1)       ����                  y�                      i(x4)       ����                  y�                      i(va_il)       ����                  y�                       	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CACsweep        XYZ[\]^_               
                       ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                      v(iv_vl)       ����                  y�                     	i(va_ix1)       ����                  y�                     i(x4)       ����                  y�                     i(va_il)       ����                  y�                      	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  �� 
 CTranSweep       vwxyz{|}               
                       ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                       v(iv_vl)       ����                  y�                      	i(va_ix1)       ����                  y�                      i(x4)       ����                  y�                      i(va_il)       ����                  y�                       	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CACdisto        qrstu               
                           ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                       v(iv_vl)       ����                  y�                      	i(va_ix1)       ����                  y�                      i(x4)       ����                  y�                      i(va_il)       ����                  y�                       	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ă        k� ����        ��������k� ����       ��������k� ����       ��������k� ����dec     ��������k� ����       ��������               
                           ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                       v(iv_vl)       ����                  y�                      	i(va_ix1)       ����                  y�                      i(x4)       ����                  y�                      i(va_il)       ����                  y�                       	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ă        k� ����        ��������k� ����       ��������k� ����       ��������k� ����dec     ��������k� ����       ��������               
                           ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                       v(iv_vl)       ����                  y�                      	i(va_ix1)       ����                  y�                      i(x4)       ����                  y�                      i(va_il)       ����                  y�                       	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ă        k� ����        ��������k� ����       ��������k� ����       ��������k� ����dec     ��������k� ����       ��������               
                           ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                       v(iv_vl)       ����                  y�                      	i(va_ix1)       ����                  y�                      i(x4)       ����                  y�                      i(va_il)       ����                  y�                       	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ă        k� ����        ��������k� ����       ��������k� ����       ��������k� ����dec     ��������k� ����       ��������               
                           ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                       v(iv_vl)       ����                  y�                      	i(va_ix1)       ����                  y�                      i(x4)       ����                  y�                      i(va_il)       ����                  y�                       	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ă        k� ����        ��������k� ����       ��������k� ����       ��������k� ����dec     ��������k� ����       ��������               
                       	    ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                       v(iv_vl)       ����                  y�                      	i(va_ix1)       ����                  y�                      i(x4)       ����                  y�                      i(va_il)       ����                  y�                       	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CACnoise        `abcdefg               
                    
    ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                      v(iv_vl)       ����                  y�                     	i(va_ix1)       ����                  y�                     i(x4)       ����                  y�                     i(va_il)       ����                  y�                      	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  J�         k�  ����        ��������k�  ����       ��������k�  ����       ��������k� ����dec     ��������k� ����       ��������k� ����       ��������k� ����  	     ��������k� ����  
     ��������              
                        ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                      v(iv_vl)       ����                  y�                     	i(va_ix1)       ����                  y�                     i(x4)       ����                  y�                     i(va_il)       ����                  y�                      	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CFourier        ~��               
         ��                   ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                      v(iv_vl)       ����                  y�                     	i(va_ix1)       ����                  y�                     i(x4)       ����                  y�                     i(va_il)       ����                  y�                      	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CACpz        	 hijklmnop               
                       ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                      v(iv_vl)       ����                  y�                     	i(va_ix1)       ����                  y�                     i(x4)       ����                  y�                     i(va_il)       ����                  y�                      	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CDCtf         HIJKL               
                       ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                      v(iv_vl)       ����                  y�                     	i(va_ix1)       ����                  y�                     i(x4)       ����                  y�                     i(va_il)       ����                  y�                      	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CDCsens         MNOPQRSTUVW               
                       ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                       v(iv_vl)       ����                  y�                      	i(va_ix1)       ����                  y�                      i(x4)       ����                  y�                      i(va_il)       ����                  y�                       	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j                  ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                      v(iv_vl)       ����                  y�                     	i(va_ix1)       ����                  y�                     i(x4)       ����                  y�                     i(va_il)       ����                  y�                      	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CShow         �              
                       ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                      v(iv_vl)       ����                  y�                     	i(va_ix1)       ����                  y�                     i(x4)       ����                  y�                     i(va_il)       ����                  y�                      	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CShowmod         �              
                       ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                      v(iv_vl)       ����                  y�                     	i(va_ix1)       ����                  y�                     i(x4)       ����                  y�                     i(va_il)       ����                  y�                      	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  �� 
 CLinearize        k�  ����        ��������               
                       ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                      v(iv_vl)       ����                  y�                     	i(va_ix1)       ����                  y�                     i(x4)       ����                  y�                     i(va_il)       ����                  y�                      	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CParamTranSweep        �������������               
                       ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                      v(iv_vl)       ����                  y�                     	i(va_ix1)       ����                  y�                     i(x4)       ����                  y�                     i(va_il)       ����                  y�                      	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  �              ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                       v(iv_vl)       ����                  y�                      	i(va_ix1)       ����                  y�                      i(x4)       ����                  y�                      i(va_il)       ����                  y�                       	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CParamACSweep        	
               
                       ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                      v(iv_vl)       ����                  y�                     	i(va_ix1)       ����                  y�                     i(x4)       ����                  y�                     i(va_il)       ����                  y�                      	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CMonteCarlo_op        ����������������������������               
                              ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                      v(iv_vl)       ����                  y�                     	i(va_ix1)       ����                  y�                     i(x4)       ����                  y�                     i(va_il)       ����                  y�                      	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CMonteCarlo_dc        ����������������������������               
                       ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                       v(iv_vl)       ����                  y�                      	i(va_ix1)       ����                  y�                      i(x4)       ����                  y�                      i(va_il)       ����                  y�                       	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CMonteCarlo_ac        ����������������������������               
                       ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                      v(iv_vl)       ����                  y�                     	i(va_ix1)       ����                  y�                     i(x4)       ����                  y�                     i(va_il)       ����                  y�                      	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CMonteCarlo_tran        ���������������������������                
                       ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                       v(iv_vl)       ����                  y�                      	i(va_ix1)       ����                  y�                      i(x4)       ����                  y�                      i(va_il)       ����                  y�                       	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CACsens                       
                              ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                       v(iv_vl)       ����                  y�                      	i(va_ix1)       ����                  y�                      i(x4)       ����                  y�                      i(va_il)       ����                  y�                       	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j  ��  CNetworkAnalysis         !"#               
                       ����            P               y�                        v(12)       ����                  y�                       v(3)       ����                  y�                       v(4)       ����                  y�                       v(5)       ����                  y�                       v(6)       ����                  y�                       v(9)       ����                  y�                       v(7)       ����                  y�                       v(8)       ����                  y�                       v(10)       ����                  y�	                       v(11)       ����                  y�
                       v(14)       ����                  y�                       v(iv_vl)       ����                  y�                      	i(va_ix1)       ����                  y�                      i(x4)       ����                  y�                      i(va_il)       ����                  y�                       	v(iv_vx1)       ����                  y�                       i(x2)       ����                  ��  � �|p�|����m�|+j  ��  � �|p�|����m�|+j                  ����            P              33�=           ��   CDigSimResTemplate                ���       ����  ����:�0�yU>20.00n���   ����                       Arial����                       Arial����                       Arial  �   �  �                                ����  ���� ������       ����  ���� ������                 �               ����  �����       200������         0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial      �       �         �     �   �  �  Circuit1                  ����  ��    ��������                                                                                     g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     ��   CPackageAliasSuperPCBStandardDIODE3      ��Eagle	DIODE.LBRDO41-7   AC  ��Orcad 	DAX2/DO41      ��	Ultiboard	L7DIO.l55DIO_DO41              A      g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     ��SuperPCBStandardDIODE3      ��Eagle	DIODE.LBRDO41-7   AC  ��Orcad 	DAX2/DO41      ��	Ultiboard	L7DIO.l55DIO_DO41              A                                                                                          g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     ��SuperPCBStandardDIODE3      ��Eagle	DIODE.LBRDO41-7   AC  ��Orcad 	DAX2/DO41      ��	Ultiboard	L7DIO.l55DIO_DO41              A      g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     ��SuperPCBStandardDIODE3      ��Eagle	DIODE.LBRDO41-7   AC  ��Orcad 	DAX2/DO41      ��	Ultiboard	L7DIO.l55DIO_DO41              A                                �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  �                _ T�� �� E .E                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                      �  �                d�         �  @                  ���                                                  �  @  6�     <   �  <     ��                                                        6�     |   �  |     ��                                                        6�     �   �  �     ��                                                        6�     �   �  �     ��                                                        f� �      �  4     ��                                                      �      �  4   �      �  4   [title]                                       f� �   D   �  t     ��                                                      �   D   �  t   �   D   �  t   [description]                                       f� `   �   h  �     ��                                                      `   �   h  �   `   �   h  �   [id]                                       f� �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       f�      �   8    ��        	                                                   �   8       �   8  Date :       �    8  �                  f� �     �  4   	 ��        
                                              �     �  4  �     �  4  [date]                                       f�       t   8    
 ��                                                            t   8         t   8   Title :       �      �                  f�    L   �   x     ��                                                         L   �   x      L   �   x   Description :       �  �  �   �                  f�    �   �   �     ��                                                         �   �   �      �   �   �   ID :       �  �  �  T                  f�    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �  L  (                      ��������������          �     	title box    Analog Misc      �?    9 
 "�     k�  ����        ��������k�  ����       ��������k�  ����       ��������k�  ����       ��������k�  ����       ��������        9                                      ����*��� ����     ,�            title                ,�            description               ,�            id               ,�            designer               ,�            date                           ����            `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                                                                                            2         �  �              � � �                   ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                          �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   
cgs 76         47 80moh5.6 ���� � mvrd nmodel             y�                      TIME� # ) time                      y�                        v(3)      v(3)    TIME                 y�                      	i(va_ix1)�   � 	i(va_ix1)    TIME                 y�    (v(7)-v(3))                   v(IV_VL)� �   v(IV_VL)    TIME                 y�                      i(va_il)  � � i(va_il)    TIME                 y�    v(5)                   	v(IV_Vx1)� �   	v(IV_Vx1)    TIME                 y�    v(iv_vx1)*i(va_ix1)                    Pin� # )  ����TIME                 y�                        v(5)      v(5)    TIME                 y�                       i(va_d2)    � i(va_d2)    TIME                 y�                       i(va_x2)� �   i(va_x2)    TIME                 y�                       i(va_x1)�   � i(va_x1)    TIME                 y�                       i(va_d1)  � @ i(va_d1)    TIME                           2         �  �           Time  � � �                   ����                       Arial����                       Arial                              ����  ����ё�[W?1.425662e-003����       ����  ����� �6lD?6.109980e-004��;]       ����  �������հ	@3.211344e+000������      ����  ������>��Nڿ-4.110512e-001������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     1m  0                            100   100                                                             1m  0                            100   100                                1m  0                            100   100                                1m  0                            100   100                                                 
                 1m  0                            100   100                            ��   CPartPackage     ��   CPackageg   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     ����   ���/� ��g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     ����   ��A
>D ��g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     ����   ���ՙ ��g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     ����      ��   CMiniPartPin    ����C+C+     PASC+�      ��   ����C-C-     PASC-�     capacitor_genericcapacitor_generic                          ��    ����11     PAS1�      ��   ����22     PAS2�     BatteryBattery                          ��    ����R+R+     PASR+      ��   ����R-R-     PASR-     RR                          ��    ����GndGnd     GNDGnd}      GndGnd                  ��    ����M+M+     PASM+i      ��   ����M-M-     PASM-j     	voltmeter	voltmeter                          ��    ����M+M+     PASM+2      ��   ����M-M-     PASM-3     Ammeter2Ammeter2                       � ��    ����D+D+     PASA       ��   ����D-D-     PASK       r   ��   CPackagePin 1 D+PAS  AA� 2 D-PAS  AKDiodeDiode	Fairchild      1n4007 D1n4007D4            diode-21n40071n4007                       � ��    ����D+D+     PASA       ��   ����D-D-     PASK       �  � 1 D+PAS  AA� 2 D-PAS  AKDiodeDiode	Fairchild      1n4007 D1n4007D3            diode-21n40071n4007                          ��    ����SW+4     PASSW+=      ��   ����SW-5     PASSW->     switch_timeswitch_time                          ��    ����SW+4     PASSW+=      ��   ����SW-5     PASSW->     switch_timeswitch_time                          ��    ����SW+4     PASSW+=      ��   ����SW-5     PASSW->     switch_timeswitch_time                          ��    ����L+L+     PASL+K      ��   ����L-L-     PASL-L     InductorInductor                          ��    ����M+M+     PASM+0      ��   ����M-M-     PASM-1     AmmeterAmmeter                          ��    ����M+M+     PASM+k      ��   ����M-M-     PASM-l     
Voltmeter2
Voltmeter2                       � ��    ����D+D+     PASA       ��   ����D-D-     PASK       w   � 1 D+PAS  AA� 2 D-PAS  AKDiodeDiode	Fairchild      1n4007 D1n4007D2            diode-21n40071n4007                       � ��    ����D+D+     PASA       ��   ����D-D-     PASK       }  � 1 D+PAS  AA� 2 D-PAS  AKDiodeDiode	Fairchild      1n4007 D1n4007D1            diode-21n40071n4007                          ��    ����M+M+     PASM+2      ��   ����M-M-     PASM-3     Ammeter2Ammeter2                          ��    ����SW+4     PASSW+=      ��   ����SW-5     PASSW->     switch_timeswitch_time                                                                                                                                                                                                           ��    �Z�P��,�                        ��                                                                                                            (f    x=f � �'f                           �(f                            ,�e    �f � ��e                           ��e                                     �  � ���� �                         .I                                                                                                       .I a    MVA_IL.I +j�6
MV                        <
                              ��    P �� �� �!�                        �"�                                             �                           �                                       h     �&   h                         �%                            �     � �� �� (�K                        �                              ��    ��������P��                        ��                            �V�    (W�`W��W��W�                        �Y�                            Їl    `�l(�l`-j �W                         �W                            t�@
    L �k��
>ENDDATA
                        
JV1                            p�<        ��<x�                           �                            \       |     ��                                                                           �rP��                                 2 2 2 2 d                                                                       