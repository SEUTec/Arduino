    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz      ��  CPart       �     �      �     �              Inductor��  CIntPin    ��  CWire     �        �
       �   �   �      �   �   �              R �   �    �   
   �       �   �   �      �   �   �              R�    �    �       6   ��   CBehPin    L-      ����L-����                        ���     R+        ����R+����                        �� 6    6  ��  CExtPin    ��  CVertex    	      ��  CSegment   �1    	  @                               �   R+  �   �    	  �   �    �7    	  �    �    �&   �  �    �   �6   �  `                  �
    �#      �   �   �+      `   $    	    #     " �   # �"   `  �   �   �)   `      (        '     &                         �"   �8   �  �   �   �*   �      ,    
    +     * �#   + �   �  �
   .                                          @  R-    	  @         RLs     ��   CPin                    ��                                                           @   R+0�                   ��                                                          �   R-��  TLine     �   �����     ��                                                        3�    �   �����     ��                                                        3�    �   �����     ��                                                        3�    x   �����     ��                                                        3�    x   ����l     ��                                                        3�    `       X     ��                                                        3�     @       X     ��                                                        3�    `   ����l    	 ��        	                                                3�     �       �    
 ��        
                                                ��  
 TTextField     t   �   �     ��                                                           t   �   �       t   �   �   [resistance]       `	  �  �	  2      `   �   �   =�     @   �   d     ��                                                           @   �   d       @   �   d   	[refname]       `	     
  �          t   $    1 2 4 5 6 7 8 9 : ; < > ?  �  resistor    resistor DINMiscellaneous      �?       ��  CResistorBehavior     ��  CValue �����������?0.1      ��������B� ���� 27     ��������B� ����       ��������B� ����       �������� R+R-  �    R-      ����R-����                        �� resistor                 G Passive   Generic   RLsRLs          ����    R ��   CPartPin    ����R+R+      PASAR+sl����H�   ����R-R-      PASAR-�sl����Passivedefault resistor, 1KGeneric              7 �   
    �       _      �      _      �              capacitor_generic�       L 3 K �    !       �  C-�  �   �-   �  �   �   �.   �  �   �   �'      �   �   T �,      �   U    	         �   T �9   `  �   �    X �	   `  �   Y             W         S     R     �   �/    	  �   �   \ �    	  `   ]             �!   �:   �  �   �	   ` �!   �  �   a    
         �$   �0   �  �   �   d �   �  `   e            c     `     _     \     [     R     Q     P                   �   C+�   �  �         C1     0�                   ��                                                           �   C-0�                   ��                                                          @   C+3�     @       �      ��    ��                                                3�     �   �����     ��                                                        3�     �   �����     ��    ��                                                3�     �       �     ��    p�H                                                =� 0   t   �   �     ��                                                       0   t   �   �   0   t   �   �   [capacitance]       0    �  �      `   �   �   =� 0   @   �   d     ��                                                       0   @   �   d   0   @   �   d   	[refname]       0  �  �             �   $    i j k l m     n       g h  �  	Capacitor     Miscellaneous      �?       ��  CCapacitorBehavior     B� '  �h㈵��>10u      ��������B� ���� x     ��������B� ����       ��������B� ����       �������� C+C- �     C+        ����C+����                        ���    C-      ����C-����                        �� 	capacitor   N           u v Passive   Generic   C1C1          ����  C H�    ����C+C+      PASAC+    ����H�   ����C-C-      PASAC-    ����Passive Generic              7 �   
   �	       �   �   �      �   �   �              resistor_generic�        z 3 y �    V        �   R+  �   %       @  R-                RCp     0�                    ��                                                           @   R+0�                   ��                                                          �   R-3�     �   �����     ��    ��                                                3�    �   �����     ��                                                        3�    �   �����     ��    ��                                                3�    x   �����     ��    p�H                                                3�    x   ����l     ��                                                       3�    `       X     ��    D�H                                                3�     @       X     ��                                                       3�    `   ����l    	 ��        	                                                3�     �       �    
 ��        
                                                =�     t   �   �     ��                                                           t   �   �       t   �   �   [resistance]       �  |  h        `   �   �   =�     @   �   d     ��                                                           @   �   d       @   �   d   	[refname]       �  �  H  �          t   $    ~  � � � � � � � � � � �  �  resistor    resistor DINMiscellaneous      �?       @�     B� ����     j�@100K      ��������B� ���� 27     ��������B� ����       ��������B� ����       �������� R+R- �     R+        ����R+����                        ���    R-      ����R-����                        �� resistor   N           � � Passive   Generic   RCpRCp          ����    R H�    ����R+R+      PASAR+    ����H�   ����R-R-      PASAR-    ����Passive Generic              7 �   
   �       _   �  �      _   �  �              
Voltmeter2�        � 3 � �    Z    `   `   M+k  �   )   `   �  M-l                 V_RLoad    
 0�                    ��                                                               M+0�                   ��                                                          �   M-3�     �       �     ��    ��                                                3�             <     ��                                                        3�    $      4     ��    ��                                                3�    ,      ,     ��    p�H                                                3�    �      �     ��               	FIXED_ROT                                        �� 
 TRectangle     <   �   �                  ����                                             <   �   �   =�    D   �   x     ��                                                         D   �   x      D   �   x   [value]         �  �  �     D   �   x   =� 8      �   0    	 ��        	                                               8      �   0   8      �   0   	[refname]       �  D  P  �  8      �   0    � � � � � � �     �       �   � 
     Voltemeter-Vert    Voltemeter-Vert_smallMiscellaneous      �?       ��   CVoltmeterBehavior     B� ����   ��l�-2.68      �������� M+M- �     M+        ����M+����                        ���    M-      ����M-����                        ��	voltmeter	voltmeter   _            � � Analog Meters   Generic   V_RLoadV_RLoad          ����  IVm H�    ����M+M+      PASAM+    ����H�   ����M-M-      PASAM-    ����Analog MetersVoltmeter-verticalGeneric              7 	 �   
   �       �   �  �      �   �  �              vcswitch�    �     �    �     �           �   �           �   �               Gnd� �    �   �      �   �   �      �          �     �   � �3          � �   �;          �   �          �         �     �   �5   �      � �   �   �  �   �         �          �     �      �     �   �%          �         �                          `       Gnd}   `             gnd1     0�                    ��                                                               Gnd3�                   ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        3�         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        3�    ,   4   ,     ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        3�    8   (   8     ��    p�Z         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         � � � �   �      Ground    
Ground DINMiscellaneous      �?       ��   CGroundBehavior       Gnd �     Gnd        ����Gnd����                        ��gndgnd                 � Analog Meters   Generic   gnd1gnd1          ����  gnd H�    ����GndGnd      GNDAGnd    ����SourcesGroundGeneric              0 � �   �    �   �����   �  �  �����   �  �              voltage_source�    �    �   �   � Ctrl �  �    3      ����3����                        ���     V+        ����V+����                        �� Ctrl   � Ctrl � �    �       �
   �   � �2      `	   �   � �4      `	   �   � �$      �
   �            �         �                           V+g  �   �       �  V-h      `	         V1     0�                   ��                                                           `   V+0�                   ��                                                          �   V-��  TEllipse     �   �����                   ����                                         �����       �   �����       �   3�    �   �����     ��    ��)                                                3�     �       �     ��    ��`                                                3�     �       �     ��    ��)                                                3�     \       �     ��    p�Z                                                3� �����   
   �    
 ��               	FIXED_ROT                                        =� \   `   \   `     ��                                                      \   `   \   `   \   `   \   `           4  �
  4  �
                =� 0   �   �   �     ��        	                                               0   �   �   �   0   �   �   �   [dc]       �    �  �          p   @   =� 0   \   �   �    	 ��        
                                               0   \   �   �   0   \   �   �   	[refname]       �  t
  0        ����t       �   � � � � � � � �       �     �  �  Voltage Source    Voltage Source DINRoot      �?       ��  CVSourceBehavior     B� ����        0      ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       �������� V+V- � �    V-      ����V-����                        ��volt_sourcevolt_source   +0            � � Sources   Generic   V1V1          ����       B�0            0      ��������B�0����      @5     ��������B�0            0     ��������B�0�  w���!�>0.3u     ��������B�0�  w���!�>0.3u     ��������B�0�8 �����>8u     ��������B�0p� �YVPh�>16.6u     ��������    B�0            0      ��������B�0����      @5     ��������B�0����     ��@10k     ��������B�0            0     ��������B�0            0     ��������    B�0            0      ��������B�0����      �?1     ��������B�0����      �?1     ��������B�0            0     ��������B�0����      �?1     ��������    B�0            0      ��������B�0����      �?1     ��������B�0            0     ��������B�0 N  �����>2u     ��������B�0'  ���ư>1u     ��������B�0'  ���ư>1u     ��������    B�  ���� 0 0      ��������                0      �������� ����       �������� ����       �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������               V H�    ����V+V+      PWR+AV+@cn����H�   ����V-V-      PWR-AV-   @����Sources Generic              0 �   �    �           �   �          �   �              Battery�    �    �       �       _   @  �      _   @  �              Ammeter2�      3 �    �   �  �   �   �   �                             `   �  M+2  �   f   `   `   M-3   @            I_Source    	 0�                    ��                                                           �   M+0�                   ��                                                              M-3�     �       �     ��                                                        3�     <             ��                                                        �� @   <   �����                  ����                                         ����<   @   �   3� ����x   ����L     ��                                                        ��  TPolygon  ������� �������  ��          @ @                                           ��  TPoint����H    ��b#�����T    
>DA#�����T    uT@ @ =� ����D   <   |     ��                                                      ����D   <   |   ����D   <   |   [value]         �    b     D   �   |   =� ��������B        ��                                                       ��������B      ��������B      	[refname]       �   �  ^  �     �����      
 '   ("	   Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       ��   CAmmeterBehavior     B� ����    �0@16.01      �������� M+M- �     M+        ����M+����                        ���    M-      ����M-����                        ��AmmeterAmmeter   V            ,-Analog Meters   Generic   I_SourceI_Source          ����  VAm H�    ����M+M+      PASAM+8�W����H�   ����M-M-      PASAM-��W����Analog MetersAmmeter-verticalGeneric              4  �     1       ����1����                        ��, 4   4 �       `       1�  �   �   `   �  2�   @             X1     0�                    ��                                                               10�                   ��                                                          �   23�             $     ��    ��)                                                3�     \       �     ��                                                        3�    8   0   8    	 ��    ��)                                                3�     H   @   H     ��    p�Z                                                3�     $   @   $     ��                                                       3�    \   0   \     ��    D�Z                                                3�               ���                                                      3�               ���   �Z	                                                =� `          $    
 ��        
                                               `          $   `          $   	[devname]        ����������������`          $   =� `   $      H     ��                                                       `   $      H   `   $      H   	[refname]       `  l  �    `   $      H    34569:;<    =>    8  7     Battery     Miscellaneous      �?    9 
 ��  CParamSubBehavior     B� ����      (@12      �������� 12 0�    2      ����2����                        ��BatteryBattery
 9 i             0BSources   Generic   X1X1          ������   CParamSubModelType��    BATTERY2.SUBCKT Xbattery 1 2
V1 1 2 DC {voltage}
.ENDS
   ��  	 CParmDefn    1battery voltage   ParamSubvoltageV                X H�    ����11      PASA10Ab����H�   ����22      PASA2�1b����SourcesBatteryGeneric              0 �   �    � 0  B� �     1       ����1����                        ���    4      ����4����                        ���   0    � 0 � � I�    �    �   �  1S  �   /   �      2T  �   �          3U  �   �       �  4V      `	        X2     0�                    ��                                                       @   �   10�                   ��                                                      @   `   20�                   ��                                                          `   30�                   ��                                                          �   43�     �       �     ��    ��                                                3�     `       �     ��                                                        3�     �       �    
 ���   ��                                                3� �����      �    	 ���   p�H                                                ܀ D   �   <   �                  ����                                         <   �   D   �   <   �   D   �   ��    �   �����               	   ����                                         �����      �   3� @   `   @   �     ��       
                                                3� 0   �   @   �     ��    D�H                                                3� @   �   @   �     ��                                                       3�    �   �����     ��  � �H        	FIXED_ROT                                        3�    �   4   �     ��                                                        =� `   �   �   �     ��                                                       `   �   �   �   `   �   �   �   	[refname]            �  �  T   �   �   �   =� �   �   @  �     ��                                                       `   `   �   �   `   `   �   �   	[devname]        ����������������T   `   �   �    PQRSYZ\      U]  ^W_`[TV    X �  vcswitch     Miscellaneous      �?   9 
 ?�    B� ����433333@4.8      ��������B� ����433333�?0.3     ��������B� ����      �?0.5     ��������B� ����    ��.A1meg     �������� 1234 J�    2      ����2����                        ��� Kvcswitchvcswitch
 9               Jf� KSwitches   Generic   X2X2          ����C���voltage controlled switch   VCSW{.subckt vcsw 1 2 3 4
S 1 2 3 4 switch
.model switch sw (vt={(Von+Voff)/2} vh={(Von-Voff)/2} ron={Ron} roff={Roff})
.ends   E�    1turnon voltage   ParamSubVon               E�    1turnoff voltage   ParamSubVoffV             E�    0on resistance   ParamSubRonOhm             E�    0off resistance   ParamSubRoffOhm               X H�    ����11      PASA1 � ����H�   ����22      PASA2NDDA����H�   ����33      PASA3    ����H�   ����44      PASA4�S����Switches Generic              7  G f� �    R-      ����R-����                        ��v �  7   7 �    b        �   R+  �   -       @  R-   �  �         RLoad     0�                    ��                                                           @   R+0�                   ��                                                          �   R-3�     �   �����     ��                                                        3�    �   �����     ��                                                        3�    �   �����     ��                                                        3�    x   �����     ��                                                       3�    x   ����l     ��    D�Z                                                3�    `       X     ��    ��d                                                3�     @       X     ��                                                        3�    `   ����l    	 ��        	                                                3�     �       �    
 ��        
                                                =�     t   �   �     ��                                                           t   �   �       t   �   �   [resistance]               �      `   �   �   =�     @   �   d     ��                                                           @   �   d       @   �   d   	[refname]          �  H             t   $    stuvwxyz{|}~ �  resistor    resistor DINMiscellaneous      �?       @�     B� ����     @�@1000      ��������B� ���� 27     ��������B� ����       ��������B� ����       �������� R+R- �     R+        ����R+����                        ��p resistor                �pPassive   Generic   RLoadRLoad          ����    R H�    ����R+R+      PASAR+    ����H�   ����R-R-      PASAR-DATA����Passivedefault resistor, 1KGeneric              3 { � M  �     L+        ����L+����                        ��-� �u �  3    3  �    ^        �   L+K  �          �  L-L    	  �         L1     0�                    ��                                                           @   L+0�                   ��                                                          �   L-��   TArc �����      �    
                                                           �����      �   �����      �       �       �           �� �����      �    	                                                           �����      �   �����      �       �       �           �� ����x      �                                                               ����x      �   ����x      �       �       x           �� ����`      x                                                               ����`      x   ����`      x       x       `           3� ����d   ����X     ��                                                        3� ����X   ����d     ��                                                        3� ����@   ����d     ��                                                        3�     @       `     ��        	                                                3�     �       �     ��        
                                                =� $   t   �   �     ��                                                       $   t   �   �   $   t   �   �   [Inductance]       l	  �  �	  �      \   �   |   =� $   @   �   d     ��                                                       $   @   �   d   $   @   �   d   	[refname]       l	  `  �	             �   $    ���  �  �  �  ���  �  �  �  � �  Inductor     Miscellaneous      �?    
   ��  CInductorBehavior     B� ��� `eG�|�>.7u      ��������B� ���� x     �������� L+L- �  Inductor  
              � Passive   Generic   L1L1          ����  L H�    ����L+L+      PASAL+    ����H�   ����L-L-      PASAL-    ����PassiveInductorGeneric                �  � � z  L �    � �   
 % ! %   & $    U       a " � Q S � � � � e ] � �  � ,  � � W [ ( Y _ * . c < ' <     � � /       � Z   �   ^            f                  � b ' # � �  T   ) - % V P R \ d  � � � � !  + X ` �    ��  CLetter    �M�s condensador y menys inductor, m�s sonidal.
Se suposa que la freq. en que Vrl seoidal coincideix amb f0.
Per tant f90 est� per sobre de la freq. senoidal, es a dir.
El condensador o la bobina encara han de ser una mica m�s grans.�  �	     �      ����Arial����                       Arial     ��   �Per C=10u, i L=.7u tenim sortida senoidal.
Si augmentem la freq. o incrementem L o C, la tensi� de sortida
disminueix en amplitud y es converteix en triangular.�  G  �  �      ����Arial����                       Arial            
 B�@ ����        ��������B�             0     ��������B� ����      @5     ��������B�  ʚ;�������?.1     ��������B�@ ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ���� true
     ��������B� ����  false     ��������               
                  B� ����        ��������B� ����       ��������B�  ����       ��������B�@ ����       ��������B�@ ����       ��������               
                  B� ����        ��������B� ����       ��������B�@ ����       ��������B�  ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������               
                 B� ����dec     ��������B� ����     @�@1k     ��������B� ����    ��.A1meg     ��������B� ����       20     ��������B� ���� true     ��������B� ���� true     ��������B� ���� true	     ��������B� ����  false
     ��������               
                 B�  ����        ��������B�  ����       ��������B�  ����       ��������B� ����dec     ��������B� ����       ��������B� ����       ��������B� ����  	     ��������B� ����  
     ��������               
                  	 B� ����        ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������               
                 B� ����        ��������B� ����       ��������B� ����       ��������B� ����dec     ��������B� ����       ��������               
                    B�             0      ��������B�  �$ hUMu/?240u     ��������B� �  H�����z>0.1u     ��������B� �  H�����z>0.1u     ��������B� ���� True     ��������B� ����  F     ��������B� ���� true     ��������B� ����  false     ��������               
                 B� ����     @�@1K      ��������B�  ����       ��������B�  ����       ��������B�  ����       ��������               
         ��              B�  ����        ��������              
                  B�  ����        ��������              
                                  
                 B�@ ����        ��������B�@ ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ���� true	     ��������B� ����  false
     ��������B� ���� true     ��������B� ����  false     ��������               
                 B� ����       5      ��������B� ����       5     ��������B� ����       5     ��������B� ����       5     ��������B� ����       ��������B� ����  	     ��������B� ����  
     ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ���� true     ��������B�@ ����       ��������B�@ ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����dec     ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ���� true     ��������B� ���� true     ��������B� ���� true     ��������B� ����  false     ��������B� ���� true     ��������B� ����  false      ��������B� ���� true!     ��������B� ����  false"     ��������               
                        B� ����       5      ��������B� ����       5     ��������B� ����       5     ��������B� ����       5     ��������B� ����       ��������B� ����  	     ��������B� ����  
     ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ���� true     ��������B�@ ����       ��������B�@ ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����dec     ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ���� true     ��������B� ���� true     ��������B� ���� true     ��������B� ����  false     ��������B� ���� true     ��������B� ����  false      ��������B� ���� true!     ��������B� ����  false"     ��������               
                 B� ����       5      ��������B� ����       5     ��������B� ����       5     ��������B� ����       5     ��������B� ����       ��������B� ����  	     ��������B� ����  
     ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ���� true     ��������B�@ ����       ��������B�@ ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����dec     ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ���� true     ��������B� ���� true     ��������B� ���� true     ��������B� ����  false     ��������B� ���� true     ��������B� ����  false      ��������B� ���� true!     ��������B� ����  false"     ��������               
                 B� ����       5      ��������B� ����       5     ��������B� ����       5     ��������B� ����       5     ��������B� ����       ��������B� ����  	     ��������B� ����  
     ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ���� true     ��������B�@ ����       ��������B�@ ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����dec     ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ���� true     ��������B� ���� true     ��������B� ���� true     ��������B� ����  false     ��������B� ���� true     ��������B� ����  false      ��������B� ���� true!     ��������B� ����  false"     ��������               
                 B�@ ����        ��������B�@ ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����decade     ��������B� ���� true     ��������B� ���� true     ��������B� ���� true     ��������B� ����  false     ��������               
                 B� ����        ��������B� ����       ��������B�@ ����       ��������B�  ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������B� ����       ��������               
                        B� ����dec     ��������B� ����     @�@1k     ��������B� ����    ��.A1meg     ��������B� ����       20     ��������B� ����        0     ��������B� ����        0     ��������B� ���� true	     ��������B� ���� true
     ��������B� ����      I@50     ��������B� ���� true     ��������B� ����  false     ��������               
                         / B� ���� x'     ��������B�     �-���q=1E-12     ��������B� @B -C��6?1E-4     ��������B� ���� x     ��������B� ���� x     ��������B� ���� x     ��������B� ���� x     ��������B� ���� x     ��������B� ���� x     ��������B� ���� x	     ��������B� ���� x!     ��������B� ����    �  500
     ��������B� ���� x     ��������B� ����    �  500     ��������B� ���� x$     ��������B� ���� x$     ��������B� ���� x%     ��������B� ���� x"     ��������B�  ���� x*     ��������B� ���� x     ��������B� ���� x     ��������B� ���� x     ��������B� ���� x&     ��������B� ���� x     ��������B� ���� x     ��������B� ���� x     ��������B� ���� x+     ��������B� ���� x,     ��������B� ���� x-     ��������B� ���� xg     ��������B� ���� xf     ��������B� ���� xd     ��������B� ���� xe     ��������B� ���� xh     ��������B� ���� xj     ��������B� ���� xi     ��������B� ���� xk     ��������B� ����    e��A1Gl     ��������B�             0�     ��������B� ����      @5�     ��������B� ����      @2.5�     ��������B� ����      �?.5�     ��������B� ����      @4.5�     ��������B� 
   ��&�.>1n�     ��������B� 
   ��&�.>1n�     ��������B� 
   ��&�.>1n�     ��������B� 
   ��&�.>1n�     ��������                 @a                Ariald         $� �|p�|����m�|+j      $� �|p�|����m�|+j                   ����                               ��  TSignal                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                     i(i_source)       ����                  ��                       i(v1)       ����                  ��                      
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CDCsweep       
 ����������               
                       ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                      i(i_source)       ����                  ��                       i(v1)       ����                  ��                       
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CACsweep        ��������               
                       ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                     i(i_source)       ����                  ��                       i(v1)       ����                  ��                      
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  �� 
 CTranSweep       ��������               
                       ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                      i(i_source)       ����                  ��                       i(v1)       ����                  ��                       
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CACdisto        �����               
                           ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                      i(i_source)       ����                  ��                       i(v1)       ����                  ��                       
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ނ        B� ����        ��������B� ����       ��������B� ����       ��������B� ����dec     ��������B� ����       ��������               
         �                 ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                      i(i_source)       ����                  ��                       i(v1)       ����                  ��                       
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ނ        B� ����        ��������B� ����       ��������B� ����       ��������B� ����dec     ��������B� ����       ��������               
         �                 ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                      i(i_source)       ����                  ��                       i(v1)       ����                  ��                       
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ނ        B� ����        ��������B� ����       ��������B� ����       ��������B� ����dec     ��������B� ����       ��������               
         �                 ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                      i(i_source)       ����                  ��                       i(v1)       ����                  ��                       
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ނ        B� ����        ��������B� ����       ��������B� ����       ��������B� ����dec     ��������B� ����       ��������               
         �                 ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                      i(i_source)       ����                  ��                       i(v1)       ����                  ��                       
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ނ        B� ����        ��������B� ����       ��������B� ����       ��������B� ����dec     ��������B� ����       ��������               
         �             	    ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                     i(i_source)       ����                  ��                       i(v1)       ����                  ��                      
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CACnoise        ��������               
                    
    ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                     i(i_source)       ����                  ��                       i(v1)       ����                  ��                      
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  .�         B�  ����        ��������B�  ����       ��������B�  ����       ��������B� ����dec     ��������B� ����       ��������B� ����       ��������B� ����  	     ��������B� ����  
     ��������              
                        ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                     i(i_source)       ����                  ��                       i(v1)       ����                  ��                      
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CFourier        ����               
         ��                   ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                     i(i_source)       ����                  ��                       i(v1)       ����                  ��                      
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CACpz        	 ���������               
                       ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                     i(i_source)       ����                  ��                       i(v1)       ����                  ��                      
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CDCtf         �����               
                       ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                     i(i_source)       ����                  ��                       i(v1)       ����                  ��                      
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CDCsens         �����������               
                       ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                      i(i_source)       ����                  ��                       i(v1)       ����                  ��                       
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j                  ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                     i(i_source)       ����                  ��                       i(v1)       ����                  ��                      
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CShow         �              
                       ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                     i(i_source)       ����                  ��                       i(v1)       ����                  ��                      
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CShowmod         �              
                       ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                     i(i_source)       ����                  ��                       i(v1)       ����                  ��                      
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  �� 
 CLinearize        B�  ����        ��������               
                       ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                     i(i_source)       ����                  ��                       i(v1)       ����                  ��                      
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CParamTranSweep        �������������               
                       ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                     i(i_source)       ����                  ��                       i(v1)       ����                  ��                      
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  �              ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                      i(i_source)       ����                  ��                       i(v1)       ����                  ��                       
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CParamACSweep        efghijklmnopq               
                       ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                     i(i_source)       ����                  ��                       i(v1)       ����                  ��                      
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CMonteCarlo_op        ����������� 	
               
                              ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                     i(i_source)       ����                  ��                       i(v1)       ����                  ��                      
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CMonteCarlo_dc         !"#$%&'()*+,               
                       ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                      i(i_source)       ����                  ��                       i(v1)       ����                  ��                       
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CMonteCarlo_ac        -./0123456789:;<=>?@ABCDEFGH               
                       ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                     i(i_source)       ����                  ��                       i(v1)       ����                  ��                      
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CMonteCarlo_tran        IJKLMNOPQRSTUVWXYZ[\]^_`abcd               
                       ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                      i(i_source)       ����                  ��                       i(v1)       ����                  ��                       
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CACsens        rstuvwxyz{|               
                              ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                      i(i_source)       ����                  ��                       i(v1)       ����                  ��                       
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CNetworkAnalysis        }~��������               
                       ����            P               ��                        v(ctrl)       ����                  ��                       v(3)       ����                  ��                       v(6)       ����                  ��                       v(4)       ����                  ��                       v(5)       ����                  ��                      i(i_source)       ����                  ��                       i(v1)       ����                  ��                       
v(v_rload)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j                  ����            P                 >           ��   CDigSimResTemplate                ���       ����  ����:�0�yU>20.00n���   ����                       Arial����                       Arial����                       Arial  �   �  �                                ����  ���� ������       ����  ���� ������                 �               ����  �����       200������         0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial      �       �         �     �   �  �  Circuit1                  ����  ��    ��������                                                                                                                                                             �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J hh?                H 1� �� L CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                      �  �                ��         �  @                  ���                                                  �  @  3�     <   �  <     ��                                                        3�     |   �  |     ��                                                        3�     �   �  �     ��                                                        3�     �   �  �     ��                                                        =� �      �  4     ��                                                      �      �  4   �      �  4   [title]                                       =� �   D   �  t     ��                                                      �   D   �  t   �   D   �  t   [description]                                       =� `   �   h  �     ��                                                      `   �   h  �   `   �   h  �   [id]                                       =� �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       =�      �   8    ��        	                                                   �   8       �   8  Date :       �    H  �                  =� �     �  4   	 ��        
                                              �     �  4  �     �  4  [date]                                       =�       t   8    
 ��                                                            t   8         t   8   Title :       �       �                  =�    L   �   x     ��                                                         L   �   x      L   �   x   Description :       �  �  �  �                  =�    �   �   �     ��                                                         �   �   �      �   �   �   ID :       �  �  �  P                  =�    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �  \  8                     �����������           �     	title box    Analog Misc      �?    9 
 ?�     B�  ����        ��������B�  ����       ��������B�  ����       ��������B�  ����       ��������B�  ����       ��������        9                                      ����C��� ����     E�            title                E�            description               E�            id               E�            designer               E�            date                           ����            `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                                                                                            2         �  �              � � �                   ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                          �   ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    
cgs 76         47 80moh5.6  ��?���mvrd nmodel ?
K3 �:� �     ��                      TIME� # ) time                      ��                        v(3)      v(3)    TIME                 ��                        v(6)      v(6)    TIME                 ��    (v(7)-v(3))                  
v(V_RLoad)� �   
v(V_RLoad)    TIME                 ��                        v(ctrl)  � � v(ctrl)    TIME                 ��                        v(7)      v(7)    TIME                 ��                      i(i_source)� �   i(i_source)    TIME                           2         �  �           Time  � � �             5
PV    ����                       Arial����                       Arial                              ����  �����z�`?2.035181e-003��G�6      ����  �����z�`?2.035181e-003��G�6      ����  ����1��{��%�-1.075922e+001������      ����  ����1��{��%�-1.075922e+001������                                                                                                                                                                                                                                                                                                                                             �  �                                              �                      �                                                                                                                                                                                                                                              1m  0                            100   100                                                             1m  0                            100   100                                1m  0                            100   100                                1m  0                            100   100                                                 
                 1m  0                            100   100                                ��   CMiniPartPin    ����L+L+     PASL+K      �   ����L-L-     PASL-L     InductorInductor                          �    ����11     PAS1�      �   ����22     PAS2�     BatteryBattery                          �    ����GndGnd     GNDGnd}      GndGnd                  �    ����R+R+     PASR+      �   ����R-R-     PASR-     RR                          �    ����M+M+     PASM+2      �   ����M-M-     PASM-3     Ammeter2Ammeter2                          �    ����11     PAS1S      �   ����22     PAS2T     �   ����33     PAS3U     �   ����44     PAS4V     vcswitchvcswitch                                         �    ����V+V+     PWR+V+g      �   ����V-V-     PWR-V-h     voltage_sourcevoltage_source                          �    ����R+R+     PASR+      �   ����R-R-     PASR-     resistor_genericresistor_generic                          �    ����R+R+     PASR+      �   ����R-R-     PASR-     RR                          �    ����C+C+     PASC+�      �   ����C-C-     PASC-�     capacitor_genericcapacitor_generic                          �    ����M+M+     PASM+k      �   ����M-M-     PASM-l     
Voltmeter2
Voltmeter2                                                                                                                                                                                                                                                                                                                                                              ,�e    �f � ��e                           ��e                                                                                                                                                                                                                                                                      
m1     8 8 mm l=100u w                        used                                                                                                            Ha    �_\PU�_\`\                        c\                            ?Q    �?Q�?Q@QXP                        �P                                                                                    2 2 2 2 d                                               