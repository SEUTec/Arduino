    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz    ��  CPart    �����   �  �  �����   �  �              voltage_source��  CIntPin    ��  CWire    �        �
   /   �   �      /   �   �                  Marker ��  CExtPin    ��  CVertex
   @  `   ��  CSegment    �6   @  �                    
        `      M     �  @          Ctrl1     ��   CPin                   ��                                                           `   M��  TLine     P       `     ��    ��                                                ��  TPolygon     ����    ����   ��                                                         ��  TPoint    0        �   @        �    P        �0   @            ��  
 TTextField    �����        ��                                                          �����         �����      	[refname]       �  1  �  �        �   ,               Marker     Miscellaneous      �?    +   ��   CMarkerBehavior     ��  CValue             0.0      �������� M ��  	 TModelPin ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �         �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               " Analog MiscV   Generic   Ctrl1Ctrl1          ����               Ctrl1  v(Ctrl1)  N ��   CPartPin    ����MM       A     ����RootmarkerGeneric              Ctrl1 �        �   /   �   �      /   �   �                  Marker% 	�    �      �   �    ( �      �   )                       `      M���� �  `          Ctrl1     �                   ��                                                           `   M�     P       `     ��     �                                                 �     ����    ����   ��                                                         �    0        �   @        �    P        �0   @            �    �����        ��                                                          �����         �����      	[refname]       �  Q  �  �        �   ,    -   + 2 ,      Marker     Miscellaneous      �?    +   �     �             0.0      �������� M !� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      3   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               5 Analog MiscV   Generic   Ctrl1Ctrl1          ����               Ctrl1  v(Ctrl1)  N #�    ����MM       A �������RootmarkerGeneric              Ctrl1 �      �       �   �  �      �   �  �              vcswitch�    �    
 �    :     �           �   �           �   �               Gnd; 	�    �   �  �   �#   �   �  `   ?          >     �"   �7   �  �   A �   �   �  �   C         B          >     �   > �,   �  �   �!   �1   �  `   G          F     E �   F �+      �   �   �2          K          J     I �   J �'   @  �   �   �-   @  `   O         N     M                                        `       Gnd}   `  �          gnd1     �                    ��                                                               Gnd�                   ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��    p�Z         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         Q R S U   T      Ground    
Ground DINMiscellaneous      �?       ��   CGroundBehavior       Gnd ��   CBehPin     Gnd        ����Gnd����                        ��gndgnd                 Y Analog Meters   Generic   gnd1gnd1          ����  gnd #�    ����GndGnd      GNDAGnd �)����SourcesGroundGeneric              0 9 �   :    �           �   �          �   �              Battery�    �    ] �    ^    �       _   @  �      _   @  �              Ammeter2_ �   �    a �    b    �       �   �        �   �                Inductorc �   �    �   f   8 6 e �    f   �       _      �      _      �              capacitor_generich �   :     i 0 	�    H       �  C-�  	�   �$   �  �   �   �5   �  @   n �   �.   �  @   �   q �!   �  �   r            �&   �       @   t        q     p     o     �   o �)   �	  @   v                 m                   �   C+�   �  �         Ce     �                   ��                                                           �   C-�                   ��                                                          @   C+�     @       �      ��    ��                                                �     �   �����     ��                                                        �     �   �����     ��    ��                                                �     �       �     ��    p�H                                                � 0   t   �   �     ��                                                       0   t   �   �   0   t   �   �   [capacitance]       0	    (
  �      `   �   �   � 0   @   �   d     ��                                                       0   @   �   d   0   @   �   d   	[refname]       0	  �  �	             �   $    z { | } ~            x y  �  	Capacitor     Miscellaneous      �?       ��  CCapacitorBehavior     � '  /W�'�>1.38u      ��������� ���� x     ��������� ����       ��������� ����       �������� C+C- X�     C+        ����C+����                        ��X�    C-      ����C-����                        �� 	capacitor    �           � � Passive   Generic   CeCe          ����  C #�    ����C+C+      PASAC+�rR����#�   ����C-C-      PASAC-    ����Passive Generic              6 �    f    �       �   �        �   �                Inductor� �   �    �   �    �       _   �         _   �                 capacitor_generic�    �    � �   �   �       �   �   �      �   �   �              R�    :     � 0 � 	�    L        @  R+  	�   �0      �   �   �/      @   � �   �&   @  @   �        �     �   � �*   @  @   �   � �4   @  �   �             �             �                  �   R-      �         RL     �                    ��                                                           �   R+�                   ��                                                          @   R-�     \      d     ��    ��)                                                � ����p      d     ��                                                        � ����p      |     ��    ��)                                                � �����      |     ��    p�Z                                                � �����      �     ��                                                       � �����       �     ��    D�Z                                                �     �       �     ��    ��d                                                � �����      �    	 ��    |�f	                                                �     \       @    
 ��    <�b
                                                �     t   �   �     ��                                                           t   �   �       t   �   �   [resistance]       `    �  �      `   �   �   �     @   �   d     ��                                                           @   �   d       @   �   d   	[refname]       `  �  �             t   $    � � � � � � � � � � � � �  �
  resistor    resistor DINMiscellaneous      �?       ��  CResistorBehavior     � ����      $@10      ��������� ���� 27     ��������� ����       ��������� ����       �������� R+R- X�     R+        ����R+����                        ��X�    R-      ����R-����                        �� resistor                � � Passive   Generic   RLRL          ����    R #�    ����R+R+      PASAR+JV1.����#�   ����R-R-      PASAR-�)����Passivedefault resistor, 1KGeneric              8 �    �    �       �   �  �      �   �  �              	voltmeter� �   :    � 0 	�    �           M+i  	�   P       �  M-j   @  �         IV_VRL    
 �                   ��                                                           `   M+�                   ��                                                          @  M-�     `       �     ��    ��                                                �     $      @    ��                                                        �    h      h     ��    ��                                                �    `      p     ��    p�H                                                �     4     4    ��               	FIXED_ROT                                        �� 
 TRectangle $   �   ����$                  ����                                         �����   $   $  � �����          ��                                                      �����        �����        [value]       �  8  �  �  (   D   �   x   � 4   `   �   �    	 ��        	                                               4   `   �   �   4   `   �   �   	[refname]       �  �  <  `         �   0    �   � � � � �   � � �       � 
 �  	voltmeter    voltmeter_smallMiscellaneous      �?       ��   CVoltmeterBehavior     � ����   ��{@ 6.62      �������� M+M- X�     M+        ����M+����                        ��X�    M-      ����M-����                        ��	voltmeter	voltmeter   _            � � Analog Meters   Generic   IV_VRLIV_VRL          ����  IVm #�    ����M+M+      PASAM+    ����#�   ����M-M-      PASAM-    ����Analog Meters Generic              8  X�     C+        ����C+����                        ��� �  8  � 8 � 	�    �#   `  @   �   � �   �  @   �                          �   C-    	�   �    �  �   C+�l� `  �         C     �                   ��                                                           @   C-�                   ��                                                      �   @   C+� �   @   `   @      ��                                                       � `   `   `         ��    p�H                                                � @   `   @         ��                                                       � @   @       @     ��    ��)                                                �     `   �   �     ��                                                           `   �   �       `   �   �   [capacitance]       `  �  �  6      `   �   �   �         �   $     ��                                                               �   $           �   $   	[refname]       `  �  �             �   $    � � � � �     �       � �    	Capacitor     Miscellaneous      �?       ��     � '  VMlS�y>0.0958u      ��������� ���� x     ��������� ����       ��������� ����       �������� C+C- � X�    C-      ����C-����                        �� 	capacitor    �           � � Passive   Generic   CC          ����  C #�    ����C+C+      PASAC+�Q����#�   ����C-C-      PASAC-h�P����Passive Generic              7 �  � X�    L-      ����L-����                        �� 7  � 7 	�    w        �   L+S  	�   �   �  �   L-�� �	  �          L     �                    ��                                                           @   L+�                   ��                                                      �   @   L-��   TArc h   ,   �   T    
                                                           h   ,   �   T   h   ,   �   T   �   @   h   @           � P   ,   h   T    	                                                           P   ,   h   T   P   ,   h   T   h   @   P   @           � 8   ,   P   T                                                               8   ,   P   T   8   ,   P   T   P   @   8   @           �     ,   8   T                                                                   ,   8   T       ,   8   T   8   @       @           � $   P      X     ��    �H                                                �    H   $   P     ��                                                        �     P   $   P     ��                                                        �     @       @     ��    ��	                                                � �   @   �   @     ��        
                                                �     \   �   |     ��                                                           \   �   |       \   �   |   [Inductance]       �	  �  (  *      \   �   |   �         �   $     ��                                                               �   $           �   $   	[refname]       �	  �  �	             �   $    � � �   �   �   �   � � �   �   �   �   �      Inductor     Miscellaneous      �?    
   ��  CInductorBehavior     � ��� ӑ�Fn4=?445.63u      ��������� ���� x     �������� L+L- X�     L+        ����L+����                        ���  Inductor  
  �           � � Passive   Generic   LL          ����  L #�    ����L+L+      PASAL+    ����#�   ����L-L-      PASAL-�,�����PassiveInductorGeneric              6  X�    2      ����2����                        ��� X�    L-      ����L-����                        ���  6  d 6 	�    �3      @   �   �"   �  @    �   �   �                     �                    �   L+K  	�   u   �  �   L-L      �          Le     �                    ��                                                           @   L+�                   ��                                                      �   @   L-� �����  �����   
                                                           h   ,   �   T   h   ,   �   T   �   @   h   @           � �����  �����   	                                                           P   ,   h   T   P   ,   h   T   h   @   P   @           � x����  �����                                                              8   ,   P   T   8   ,   P   T   P   @   8   @           � `����  x����                                                                  ,   8   T       ,   8   T   8   @       @           � $   P      X     ��    ��                                                �    H   $   P     ��                                                        �     P   $   P     ��    ��                                                �     @       @     ��    p�H	                                                � �   @   �   @     ��       
                                                �     \   �   |     ��                                                           \   �   |       \   �   |   [Inductance]          �    *      \   �   |   �         �   $     ��                                                               �   $           �   $   	[refname]          �  �             �   $              
  	         Inductor     Miscellaneous      �?    
   ��     � ��� �5��B��>25.4u      ��������� ���� x     �������� L+L- X�     L+        ����L+����                        ���  Inductor  
  �           � Passive   Generic   LeLe          ����  L #�    ����L+L+      PASAL+��N����#�   ����L-L-      PASAL-    ����PassiveInductorGeneric              5  X�    M-      ����M-����                        �� 5  ` 5 	�    �   �  �   �$   �   �  `                          `   �  M+2  	�     `   `   M-3   @  �         VA_Ix1    	 �                    ��                                                           �   M+�                   ��                                                              M-�     �       �     ��                                                        �     <             ��                                                        À @   <   �����                  ����                                         ����<   @   �   � ����x   ����L     ��                                                        �  ������� �������  ��          @ @                                           �����H    ��b�����T    
>DA�����T    uT@ @ � ����D   <   |     ��                                                      ����D   <   |   ����D   <   |   [value]         �  �  "     D   �   |   � ��������O        ��                                                       ��������O      ��������O      	[refname]       �   �  =  ?     �����      
  !"(  #)$	   Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       ��   CAmmeterBehavior     � ����   `j	�-3.18      �������� M+M- X�     M+        ����M+����                        ��AmmeterAmmeter   V            -Analog Meters   Generic   VA_Ix1VA_Ix1          ����  VAm #�    ����M+M+      PASAM+��W����#�   ����M-M-      PASAM-8�W����Analog MetersAmmeter-verticalGeneric              4  X�     1       ����1����                        ��- 4   \ 4 [ 	�       `       1�  	�   D   `   �  2�   @  `          X1     �                    ��                                                               1�                   ��                                                          �   2�             $     ��    ��)                                                �     \       �     ��                                                        �    8   0   8    	 ��    ��)                                                �     H   @   H     ��    p�Z                                                �     $   @   $     ��                                                       �    \   0   \     ��    D�Z                                                �               ���                                                      �               ���   �Z	                                                � `          $    
 ��        
                                               `          $   `          $   	[devname]        ����������������`          $   � `   $      H     ��                                                       `   $      H   `   $      H   	[refname]       `  �  �  l  `   $      H    34569:;<    =>    8  7     Battery     Miscellaneous      �?    9 
 ��  CParamSubBehavior     � ����      (@12      �������� 12 0X�    2      ����2����                        ��BatteryBattery
 9 i             0BSources   Generic   X1X1          ������   CParamSubModelType��    BATTERY2.SUBCKT Xbattery 1 2
V1 1 2 DC {voltage}
.ENDS
   ��  	 CParmDefn    1battery voltage   ParamSubvoltageV                X #�    ����11      PASA1�1b����#�   ����22      PASA20Ab����SourcesBatteryGeneric              0 j � � �    :     �	           �   �           �   �               GndI	�    �      `            	        `       Gnd}   �  `          gnd3     �                    ��                                                               Gnd�                   ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         MNOQ  P     Ground    
Ground DINMiscellaneous      �?       V�       Gnd X�     Gnd        ����Gnd����                        ��gndgnd                 SAnalog Meters   Generic   gnd3gnd3          ����  gnd #�    ����GndGnd      GNDAGnd    ����SourcesGroundGeneric              0 �   :    8 0 �    :     �           �   �           �   �               GndV	�    �   @  �   �%   �   @  @   Z         Y                `       Gnd}   �  �          gnd4     �                    ��                                                               Gnd�                   ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��    D�H         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��    x�W         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��    X��         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         \]^`  _     Ground    
Ground DINMiscellaneous      �?       V�       Gnd X�     Gnd        ����Gnd����                        ��gndgnd                 bAnalog Meters   Generic   gnd4gnd4          ����  gnd #�    ����GndGnd      GNDAGnd    ����SourcesGroundGeneric              0 �   :     0 
 X�    V-      ����V-����                        ��BY X�     1       ����1����                        ��X�    4      ����4����                        ��Sb� � �   0    8 0 g 7 U	�    @    �   �  1S  	�   s   �      2T  	�   *          3U  	�   L      �  4V      �        X2     �                    ��                                                       @   �   1�                   ��                                                      @   `   2�                   ��                                                          `   3�                   ��                                                          �   4�     �       �     ��    ��                                                �     `       �     ��                                                        �     �       �    
 ���   ��                                                � �����      �    	 ���   p�H                                                ��  TEllipse D   �   <   �                  ����                                         <   �   D   �   <   �   D   �   À    �   �����               	   ����                                         �����      �   � @   `   @   �     ��       
                                                � 0   �   @   �     ��    D�H                                                � @   �   @   �     ��                                                       �    �   �����     ��  � �H        	FIXED_ROT                                        �    �   4   �     ��                                                        � T   �   �   �     ��                                                       T   �   �   �   T   �   �   �   	[refname]       �  |  l        (   t   L   �     �  <    ��                                                       T   `   �   �   T   `   �   �   	[devname]        ����������������       �   (    lmnovwy      qz  {s|}xpr    u �  vcswitch     Miscellaneous      �?   9 
 ?�    � ����������@4.9      ��������� �����������?1.1     ��������� ����      �?0.5     ��������� ����    ��.A1meg     �������� 1234 f� X�    3      ����3����                        ��gvcswitchvcswitch
 9               f� �gSwitches   Generic   X3X3          ����C���voltage controlled switch   VCSW{.subckt vcsw 1 2 3 4
S 1 2 3 4 switch
.model switch sw (vt={(Von+Voff)/2} vh={(Von-Voff)/2} ron={Ron} roff={Roff})
.ends   E�    1turnon voltage   ParamSubVon               E�    1turnoff voltage   ParamSubVoffV             E�    0on resistance   ParamSubRonOhm             E�    0off resistance   ParamSubRoffOhm               X #�    ����11      PASA1�A�����#�   ����22      PASA2    ����#�   ����33      PASA3�����#�   ����44      PASA48 � ����Switches Generic              Ctrl1   X�     V+        ����V+����                        ���" 5  Ctrl1    Ctrl1 d	�               V+g  	�   [      �  V-h   @  �         V1     �                   ��                                                           `   V+�                   ��                                                          �   V-t�     �   �����                   ����                                         �����       �   �����       �   �    �   �����     ��    ��)                                                �     �       �     ��    ��`                                                �     �       �     ��    ��)                                                �     \       �     ��    p�Z                                                � �����   
   �    
 ��               	FIXED_ROT                                        � \   `   \   `     ��                                                      \   `   \   `   \   `   \   `           T  �  T  �                � 0   �   �   �     ��        	                                               0   �   �   �   0   �   �   �   [dc]       �  P    �          p   @   � 0   \   �   �    	 ��        
                                               0   \   �   �   0   \   �   �   	[refname]       �  �  P  T      ����t       �  ��������      �    � �  Voltage Source    Voltage Source DINRoot      �?       ��  CVSourceBehavior     � ����        0      ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       �������� V+V- �evolt_sourcevolt_source   +0            �eSources   Generic   V1V1          ����       �0            0      ���������0����      @5     ���������0            0     ���������0�  H�����z>0.1u     ���������0�  H�����z>0.1u     ���������0@ �h㈵��>20u     ���������0� �h㈵�?40u     ��������    �0            0      ���������0����      @5     ���������0����     ��@10k     ���������0            0     ���������0            0     ��������    �0            0      ���������0����      �?1     ���������0����      �?1     ���������0            0     ���������0����      �?1     ��������    �0            0      ���������0����      �?1     ���������0            0     ���������0 N  �����>2u     ���������0'  ���ư>1u     ���������0'  ���ư>1u     ��������    �  ���� 0 0      ��������                0      �������� ����       �������� ����       �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������               V #�    ����V+V+      PWR+AV+ � ����#�   ����V-V-      PWR-AV-NDDA����Sources Generic                \   <   ` 8   J W  &       � � � �     d i    :  ^ b f � � '  '                             M O � � I K � � �  p E r v  n C ) G A ? Zt 8 # 8   D Y@         >      (         [      *           L� u s � m   � N   w � J F P q � � H L � � o  B    ��  CLetter    OLC formen un filtro per obtenir tensi� senoidal a la RL.
fr=1/(2*pi*sqrt(L*C))�  G
    '    �?����Arial����                       Arial     Á   Ctrl1�     z  �      ����Arial����                       Arial     Á   0�  �  �  k    �?����Arial����                       Arial     Á   4�  p  E  �    �?����Arial����                       Arial     Á   0`  (  �  �    �?����Arial����                       Arial     Á   5�  �  E  +    �?����Arial����                       Arial     Á   6     e  �    �?����Arial����                       Arial     Á   Ctrl1P     :  �    �?����Arial����                       Arial     Á   0P  �  �  [    �?����Arial����                       Arial     Á	   7�  �  �  S    �?����Arial����                       Arial     Á
   8�  �    S    �?����Arial����                       Arial            
 �@ ����        ���������             0     ��������� ����      @5     ���������  ʚ;�������?.1     ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ���� true
     ��������� ����  false     ��������               
                  � ����        ��������� ����       ���������  ����       ���������@ ����       ���������@ ����       ��������               
                  � ����        ��������� ����       ���������@ ����       ���������  ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������               
                 � ����dec     ��������� ����     @�@1k     ��������� ����    ��.A1meg     ��������� ����       20     ��������� ���� true     ��������� ���� true     ��������� ���� true	     ��������� ����  false
     ��������               
                 �  ����        ���������  ����       ���������  ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����  	     ��������� ����  
     ��������               
                  	 � ����        ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������               
                 � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                    �             0      ���������  >I hUMu??480u     ��������� �  H�����z>0.1u     ��������� �  H�����z>0.1u     ��������� ���� True     ��������� ����  F     ��������� ���� true     ��������� ����  false     ��������               
                 � ����     @�@1K      ���������  ����       ���������  ����       ���������  ����       ��������               
         ��              �  ����        ��������              
                  �  ����        ��������              
                                  
                 �@ ����        ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ���� true	     ��������� ����  false
     ��������� ���� true     ��������� ����  false     ��������               
                 � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                        � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                 � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                 � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                 �@ ����        ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����decade     ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������               
                 � ����        ��������� ����       ���������@ ����       ���������  ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������               
                        � ����dec     ��������� ����     @�@1k     ��������� ����    ��.A1meg     ��������� ����       20     ��������� ����        0     ��������� ����        0     ��������� ���� true	     ��������� ���� true
     ��������� ����      I@50     ��������� ���� true     ��������� ����  false     ��������               
                         / � ���� x'     ���������     �-���q=1E-12     ��������� @B -C��6?1E-4     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x	     ��������� ���� x!     ��������� ����    �  500
     ��������� ���� x     ��������� ����    �  500     ��������� ���� x$     ��������� ���� x$     ��������� ���� x%     ��������� ���� x"     ���������  ���� x*     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x&     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x+     ��������� ���� x,     ��������� ���� x-     ��������� ���� xg     ��������� ���� xf     ��������� ���� xd     ��������� ���� xe     ��������� ���� xh     ��������� ���� xj     ��������� ���� xi     ��������� ���� xk     ��������� ����    e��A1Gl     ���������             0�     ��������� ����      @5�     ��������� ����      @2.5�     ��������� ����      �?.5�     ��������� ����      @4.5�     ��������� 
   ��&�.>1n�     ��������� 
   ��&�.>1n�     ��������� 
   ��&�.>1n�     ��������� 
   ��&�.>1n�     ��������                 @~                Ariald         � �|p�|����m�|+j      � �|p�|����m�|+j                   ����                             	 ��  TSignal                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                     	i(va_ix1)       ����                  �                      	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CDCsweep       
 ����������               
                       ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                      	i(va_ix1)       ����                  �                       	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CACsweep        ��������               
                       ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                     	i(va_ix1)       ����                  �                      	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  �� 
 CTranSweep       	
               
                       ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                      	i(va_ix1)       ����                  �                       	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CACdisto                       
                           ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                      	i(va_ix1)       ����                  �                       	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  �        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                           ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                      	i(va_ix1)       ����                  �                       	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  �        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                           ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                      	i(va_ix1)       ����                  �                       	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  �        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                           ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                      	i(va_ix1)       ����                  �                       	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  �        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                           ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                      	i(va_ix1)       ����                  �                       	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  �        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                       	    ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                     	i(va_ix1)       ����                  �                      	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CACnoise        ��������               
                    
    ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                     	i(va_ix1)       ����                  �                      	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  e�         �  ����        ���������  ����       ���������  ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����  	     ��������� ����  
     ��������              
                        ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                     	i(va_ix1)       ����                  �                      	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CFourier                       
         ��                   ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                     	i(va_ix1)       ����                  �                      	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CACpz        	 �������                
                       ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                     	i(va_ix1)       ����                  �                      	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CDCtf         �����               
                       ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                     	i(va_ix1)       ����                  �                      	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CDCsens         �����������               
                       ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                      	i(va_ix1)       ����                  �                       	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j                  ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                     	i(va_ix1)       ����                  �                      	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CShow                       
                       ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                     	i(va_ix1)       ����                  �                      	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CShowmod                       
                       ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                     	i(va_ix1)       ����                  �                      	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  �� 
 CLinearize        �  ����        ��������               
                       ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                     	i(va_ix1)       ����                  �                      	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CParamTranSweep         !               
                       ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                     	i(va_ix1)       ����                  �                      	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  �              ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                      	i(va_ix1)       ����                  �                       	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CParamACSweep        �������������               
                       ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                     	i(va_ix1)       ����                  �                      	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CMonteCarlo_op        "#$%&'()*+,-./0123456789:;<=               
                              ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                     	i(va_ix1)       ����                  �                      	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CMonteCarlo_dc        >?@ABCDEFGHIJKLMNOPQRSTUVWXY               
                       ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                      	i(va_ix1)       ����                  �                       	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CMonteCarlo_ac        Z[\]^_`abcdefghijklmnopqrstu               
                       ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                     	i(va_ix1)       ����                  �                      	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CMonteCarlo_tran        vwxyz{|}~������������������               
                       ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                      	i(va_ix1)       ����                  �                       	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CACsens        �����������               
                              ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                      	i(va_ix1)       ����                  �                       	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j  ��  CNetworkAnalysis        �����������               
                       ����            P              	 �                        v(ctrl1)       ����                  �                       v(4)       ����                  �                       v(5)       ����                  �                       v(6)       ����                  �                       v(7)       ����                  �                       v(8)       ����                  �                       i(v1)       ����                  �                      	i(va_ix1)       ����                  �                       	v(iv_vrl)       ����                      � �|p�|����m�|+j      � �|p�|����m�|+j                  ����            P                 >          ��   CDigSimResTemplate                ���       ����  ����:�0�yU>20.00n���   ����                       Arial����                       Arial����                       Arial  �   �  �                                ����  ���� ������       ����  ���� ������                 �               ����  �����       200������         0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial      �       �         �     �   �  �  Circuit1                  ����  ��    ��������                                                                                                                                                                                                             �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            N  M�                H 1� �� L AE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                      �  �                À         �  @                  ���                                                  �  @  �     <   �  <     ��                                                        �     |   �  |     ��                                                        �     �   �  �     ��                                                        �     �   �  �     ��                                                        � �      �  4     ��                                                      �      �  4   �      �  4   [title]                                       � �   D   �  t     ��                                                      �   D   �  t   �   D   �  t   [description]                                       � `   �   h  �     ��                                                      `   �   h  �   `   �   h  �   [id]                                       � �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       �      �   8    ��        	                                                   �   8       �   8  Date :       �    H  �                  � �     �  4   	 ��        
                                              �     �  4  �     �  4  [date]                                       �       t   8    
 ��                                                            t   8         t   8   Title :       �       �                  �    L   �   x     ��                                                         L   �   x      L   �   x   Description :       �  �  �  �                  �    �   �   �     ��                                                         �   �   �      �   �   �   ID :       �  �  �  P                  �    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �  \  8                     >?@ABCDEFHIJKL          G     	title box    Analog Misc      �?    9 
 ?�     �  ����        ���������  ����       ���������  ����       ���������  ����       ���������  ����       ��������        9                                      ����C��� ����     E�            title                E�            description               E�            id               E�            designer               E�            date                           ����            `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                                                                                            2         �  �              � � �                   ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                            �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                   
cgs 76         47 80moh5.6 >ENDDATAmvrd nmodel 12000000-0     �                      TIME� # ) time                      �                        i(v1)� < � i(v1)    TIME                 �                       	i(va_ix1)�   � 	i(va_ix1)    TIME                 �                        v(ctrl1)      v(ctrl1)    TIME                 �                        v(6)      v(6)    TIME                 �    (v(6)-v(3))                  	v(IV_VRL)� �   	v(IV_VRL)    TIME                           2         �  �           Time  � � �           JV1.    ����                       Arial����                       Arial                              ����  �����z�`?2.035181e-003��G�6      ����  �����z�`?2.035181e-003��G�6      ����  ����1��{��%�-1.075922e+001������      ����  ����1��{��%�-1.075922e+001������                                                                           �                      �                                                                                                                                                                          �  �                                                                                                                                                                                                                                                                                                                  �  �                                                                                                                          1m  0                            100   100                                                             1m  0                            100   100                                1m  0                            100   100                                1m  0                            100   100                                                 
                 1m  0                            100   100                                ��   CMiniPartPin    ����V+V+     PWR+V+g      a�   ����V-V-     PWR-V-h     voltage_sourcevoltage_source               �  �     a�    ����11     PAS1�      a�   ����22     PAS2�     BatteryBattery               �  �     a�    ����GndGnd     GNDGnd}      GndGnd                  a�    ����M+M+     PASM+2      a�   ����M-M-     PASM-3     Ammeter2Ammeter2                   �     a�    ����11     PAS1S      a�   ����22     PAS2T     a�   ����33     PAS3U     a�   ����44     PAS4V     vcswitchvcswitch                           �  �  �     a�    ����GndGnd     GNDGnd}      GndGnd                  a�    ����MM       ��������MarkerMarker                  a�    ����GndGnd     GNDGnd}      GndGnd                  a�    ����MM       ��������MarkerMarker                  a�    ����C+C+     PASC+�      a�   ����C-C-     PASC-�     capacitor_genericcapacitor_generic               �  �     a�    ����L+L+     PASL+K      a�   ����L-L-     PASL-L     InductorInductor                          a�    ����R+R+     PASR+      a�   ����R-R-     PASR-     RR                          a�    ����M+M+     PASM+i      a�   ����M-M-     PASM-j     	voltmeter	voltmeter                          a�    ����L+L+     PASL+K      a�   ����L-L-     PASL-L     InductorInductor                          a�    ����C+C+     PASC+�      a�   ����C-C-     PASC-�     capacitor_genericcapacitor_generic                                                             Ctrl1�                   0�                   41                   02                   5                   6i                   Ctrl1j                   0k                   7�                    8�                                                                                                                              
m1     8 8 mm l=100u w                        used                                                                                                            ,�e    �f � ��e                           ��e                                                                                                                                                                                                                                                                                                                                                                                                                                      h�    ���������                        ��                            ���    p�������                        q�                            �2�    �Q�R�XR��R�                        T�                            (f    x=f � �'f                           �(f                                     �  � ���� �                         .I                              �N    xW�WX�p 4M                        ЮW                                                                                    2 2 2 2 d                                                       