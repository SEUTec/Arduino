    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz    ��  CPart    �����   �  �  �����   �  �              voltage_source��  CIntPin    ��  CWire    �        �   /   �   �      /   �   �                  Marker ��  CExtPin    ��  CVertex    
   
   ��  CSegment
    �    
  �
                          `      M     �	   	          VControl     ��   CPin                   ��                                                           `   M��  TLine     P       `     ��    ���                                                 ��  TPolygon     ����    ����   ��                                                         ��  TPoint    0    Amm�   @        �    P        �0   @    P�X    ��  
 TTextField       �   ,     ��                                                             �   ,         �   ,   	[refname]       �	  	  s  �	        �   ,               Marker     Miscellaneous      �?    +   ��   CMarkerBehavior     ��  CValue             0.0      �������� M ��  	 TModelPin ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �         �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               " Analog MiscV   Generic   VControlVControl          ����               VControl  v(VControl)  N ��   CPartPin    ����MM       A  ������RootmarkerGeneric              VControl �        �   /   �   �      /   �   �                  Marker% 	�    �3       
   �)   ( �2      �
   )                       `      M     �   	          VControl     �                   ��                                                           `   M�     P       `     ��    ���                                                 �     ����    ����   ��                                                         �    0        �   @    ����    P    H���0   @    ��    �       �   )     ��                                                             �   )         �   )   	[refname]       �  	  t  �	        �   ,    -   + 2 ,      Marker     Miscellaneous      �?    +   �     �             0.0      �������� M !� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      3   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               5 Analog MiscV   Generic   VControlVControl          ����               VControl  v(VControl)  N #�    ����MM       A Teu ����RootmarkerGeneric              VControl �        �	   /   �   �      /   �   �                  Marker7 	�    �4   �  `	   �   : �   �   
   ;                 	        `      M     `  @          VControl     �                   ��                                                           `   M�     P       `     ��    ���                                                 �     ����    ����   ��                                                         �    0      �   @      �    P        �0   @            �       �   ,     ��                                                             �   ,         �   ,   	[refname]       x  X    	        �   ,    ?   = D >      Marker     Miscellaneous      �?    +   �     �             0.0      �������� M !� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      E   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               G Analog MiscV   Generic   VControlVControl          ����               VControl  v(VControl)  N #�    ����MM       A     ����RootmarkerGeneric              VControl  �      �       �   �  �      �   �  �              vcswitch�    �     �    L     �           �   �           �   �               GndM 	�    �$          �#   �0   @      Q �/   �   @      S          R          P     �!   P �&   `      �   �(    
      W �   X �+   �
      Y �   �   �
      [         Z              �   �    
      ]         X          V     U �   �   `  `   _          V              �    �.          a         P                 `       Gnd}   �             gnd1     �                    ��                                                               Gnd�                   ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��    ���          AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��    ���          AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��    ��K         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         c d e g   f      Ground    
Ground DINMiscellaneous      �?       ��   CGroundBehavior       Gnd ��   CBehPin     Gnd        ����Gnd����                        ��gndgnd                 k Analog Meters   Generic   gnd1gnd1          ����  gnd #�    ����GndGnd      GNDAGnd    ����SourcesGroundGeneric              0 K �   L    �       �   �  �      �   �  �              vcswitch�    �    o �   p   �       �   �         �   �                 1n4007�    �	    �   t  	 �       _   @  �      _   @  �              Ammeter2�    �    �   x   �       �   �  �      �   �  �              	voltmeter�    �    { �    |    �       S   �  ,      S   �  ,              Ammeter} �   �
    �    �   
 �       �   �  �       �   �  �               resistor_generic� �   x   � 4 	�    �!   �  @   �	   �   �  @   �  
      �      
              �   R+    	�   �    @  @   �   � �   �
  @   �   �,   �
  �   �"   �:   �	  �   �        �     �'   � �*   �
  �   �   �   �
  `   �         �     �   �-   `	  �   �        �     �         �     �     �+   �7   �
      � �   �#   �      �        �         �     �                  �  �   R-    �  �          RL     �                    ��                                                           @   R+�                   ��                                                      �   @   R-� d   @   \   P     ��    ���                                                 � P   0   \   P     ��                                                        � P   0   D   P     ��    ���                                                 � 8   0   D   P     ��    (�K                                                � 8   0   ,   P     ��                                                       �     0      @     ��    ��K                                                �     @      @     ��                                                       �     0   ,   P    	 ��        	                                                � d   @   �   @    
 ��        
                                                �     `   �   �     ��                                                           `   �   �       `   �   �   [resistance]       �  �  �  .      `   �   �   �         t   $     ��                                                               t   $           t   $   	[refname]       �  �  I  +          t   $    � � � � � � � � � � � � �      resistor    resistor DINMiscellaneous      �?       ��  CResistorBehavior     � ����    �ׇA50meg      ��������� ���� 27     ��������� ����       ��������� ����       �������� R+R- j� �,  R+        
  R+����                        ��j� �,  R-      
  R-����                        �� resistor   W           � � Passive   Generic   RLRL          ����    R #�    ����R+R+      PASAR+�:�    #�   ����R-R-      PASAR- �    Passive Generic              13   � j� �  M-      R  M-����                        ��
 13 
 ~ 13 	�    �	      @   �   � �   @  @   �*   �/   @      � �   � �%   @      �                 �     � �,   � �5   @  �   �$   � �1   `  �   �    
        � �   � �"   @  �   � �&   �   @  `   �         �     �   � �   �  �   � �   � �)   �  �   �                                                            �   M+    	�   �   �  �   M-       �          IRL    	 �                   ��                                                           @   M+�                   ��                                                      �   @   M-� �   @   �   @     ��    ���                                                 �     @       @     ��                                                        � 4   X   `   X     ��    ���                                                 �� 
 TRectangle        �   d                   ����                                                �   d   � ����������������  ��          @ @                                           �d   X        �X   P        �X   `        @ @ � $   $   �   L     ��                                                      $   $   �   L   $   $   �   L   [value]       l  �  Q  z  $   $   �   L   �     �����        ��                                                           �����          �����      	[refname]       `  \          �����       �   � � �   �   � � �   � 	     Ammeter    Ammeter_smallMiscellaneous      �?       ��   CAmmeterBehavior     � �t      ��> 2.99u      �������� M+M- j� �  M+        R  M+����                        ��� AmmeterAmmeter   �            � � Analog Meters   Generic   IRLIRL          ����  VAm #�    ����M+M+      PASAM+��Q    #�   ����M-M-      PASAM-��    Analog MetersAmmeterGeneric              3 �   |   �
       �   �        �   �                Inductor�    �    �    �    �   /   �      �   /   �      �               Marker� 	�    �
   `  @   �-   �8   `  �   �%   �9   @  �   �    
     �     �   � �;   �  �   �             �     �     �(   � �   `  �   �                        `      M                  VSource     �                   ��                                                           `   M� 0   `       `     ��    ���                                                 �     `       `      ��                                                         �P   `       ��@   P    ȭW�0   `    h�V�@   p          � `   P      t     ��                                                       `   P      t   `   P      t   	[refname]            �  �        �   ,    �   � � �  �  Marker     Miscellaneous      �?    +   �     �             0.0      �������� M !� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  + �             � Analog MiscV   Generic   VSourceVSource          ����               VSource  
v(VSource)  N #�    ����MM       A   ����RootmarkerGeneric              VSource � �    �    �       �   �        �   �                Inductor� �   x   � 4 	�    �        �   L+K  	�   �   �  �   L-L   �             L1     �                    ��                                                           @   L+�                   ��                                                      �   @   L-��   TArc ����,   ���T   
                                                           h   ,   �   T   h   ,   �   T   �   @   h   @           �� ����,  ����T   	                                                           P   ,   h   T   P   ,   h   T   h   @   P   @           �� ����,  ����T                                                              8   ,   P   T   8   ,   P   T   P   @   8   @           �� ����,  ����T                                                                  ,   8   T       ,   8   T   8   @       @           � $   P      X     ��    ���                                                 �    H   $   P     ��                                                        �     P   $   P     ��    ���                                                 �     @       @     ��    (�K	                                                � �   @   �   @     ��       
                                                �     \   �   |     ��                                                           \   �   |       \   �   |   [Inductance]       �    R  �      \   �   |   �         �   $     ��                                                               �   $           �   $   	[refname]       �     R  �          �   $    � �                �   �      Inductor     Miscellaneous      �?    
   ��  CInductorBehavior     � ��� {�G�zt?5m      ��������� ���� x     �������� L+L- j�     L+        ����L+����                        ��j�    L-      ����L-����                        �� Inductor  
 �           Passive   Generic   L1L1          ����  L #�    ����L+L+      PASAL+    ����#�   ����L-L-      PASAL-    ����PassiveInductorGeneric              VSource �    �    �           �   �          �   �              Battery�   �    �     �       _   @  �      _   @  �              Ammeter2�    L     0 	�    `    `   �  M+2  	�   �   `  �
   �   �   `   
                       `   `   M-3      �
         ISource    	 �                    ��                                                           �   M+�                   ��                                                              M-�     �       �     ��                                                        �     <             ��                                                        ̀ @   <   �����                  ����                                         ����<   @   �   � ����x   ����L     ��                                                        �  ������� �������  ��          @ @                                           �����H    ��b�����T    
>DA�����T    uT@ @ � ����D   <   |     ��                                                      ����D   <   |   ����D   <   |   [value]       �  L  �  �     D   �   |   � ��������B        ��                                                       ��������B      ��������B      	[refname]       �  b
  �       �����      
  !'  "(#	   Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       Ԁ     � �w��    �Rd�-2.48m      �������� M+M- j�     M+        ����M+����                        ��j�    M-      ����M-����                        ��AmmeterAmmeter   V            +,Analog Meters   Generic   ISourceISource          ����  VAm #�    ����M+M+      PASAM+   @����#�   ����M-M-      PASAM-��W����Analog MetersAmmeter-verticalGeneric              6  j�    2      ����2����                        ��, 6  6 	�    �    `       1�  	�     `   �  2�      �          X1     �                    ��                                                               1�                   ��                                                          �   2�             $     ��    ��)                                                �     \       �     ��                                                        �    8   0   8    	 ��    ��)                                                �     H   @   H     ��    p�Z                                                �     $   @   $     ��                                                       �    \   0   \     ��    D�Z                                                �               ���                                                      �               ���   �Z	                                                � `          $    
 ��        
                                               `          $   `          $   	[devname]        ����������������`          $   � `   $      H     ��                                                       `   $      H   `   $      H   	[refname]          	  �  �	  `   $      H    234589:;    <=    7  6     Battery     Miscellaneous      �?    9 
 ��  CParamSubBehavior     � ����      (@12      �������� 12 j�     1       ����1����                        ��/BatteryBattery
 9 i             A/Sources   Generic   X1X1          ������   CParamSubModelType��    BATTERY2.SUBCKT Xbattery 1 2
V1 1 2 DC {voltage}
.ENDS
   ��  	 CParmDefn    1battery voltage   ParamSubvoltageV                X #�    ����11      PASA10Ab����#�   ����22      PASA2�1b����SourcesBatteryGeneric              VSource  Aj�     L+        ����L+����                        ���  VSource   � VSource � 	�    �    �  �   L+K  	�   �       �   L-L   `            L2     �                    ��                                                       �   @   L+�                   ��                                                          @   L-�� ,����  T����   
                                                               ,   8   T       ,   8   T       @   8   @           �� ,���p  T����   	                                                           8   ,   P   T   8   ,   P   T   8   @   P   @           �� ,���X  T���p                                                              P   ,   h   T   P   ,   h   T   P   @   h   @           �� ,���@  T���X                                                              h   ,   �   T   h   ,   �   T   h   @   �   @           � |   0   �   (     ��    t                                                � �   8   |   0     ��     "                                                 � �   0   |   0     ��                                                        � �   @   �   @     ��    ���	                                                �     @   ����@     ��    ����
                                                �     \   �   |     ��                                                           \   �   |       \   �   |   [Inductance]       `    �  �      \   �   |   �         �   $     ��                                                               �   $           �   $   	[refname]       `     �  �          �   $    KLU  T  S  R  QVW  P  O  N  M   Inductor     Miscellaneous      �?    
   	�     � ��� {�G�zt?5m      ��������� ���� x     �������� L+L- Hj�    L-      ����L-����                        �� Inductor  
 �           H[Passive   Generic   L2L2          ����  L #�    ����L+L+      PASAL+    ����#�   ����L-L-      PASAL-    ����PassiveInductorGeneric              3 �    |    �       _   @  �      _   @  �              Ammeter2^�   �    `�    a   �       �   �         �   �                 1n4007b�   �    �   e  J 7 d j�    2      ����2����                        ��j�    D-      ����D-����                        �� 7  c7 	�    �   @  �                          D+   	�   �   @   	   �.   l�   @  �
   m                        @  D-    @  �         D1     �                   ��                                                           `   D+�                   ��                                                          �   D-�     �       �      ��    ���                                                 �     �   �����     ��                                                        �     �   �����     ��    ���                                                 �     `       �     ��                                                       �    �       �     ��    ��K                                                �     �   �����     ��    ��K                                                �     �       �     ��    JL1.                                                � 0   `   �   �    	 ��        	                                               0   `   �   �   0   `   �   �   	[devname]        �������������������������      � -   �   �   �    
 ��        
                                               -   �   �   �   -   �   �   �   	[refname]       �  [  P  	  ����   �   <    qrstuvw    xy          op �  diode     Miscellaneous      �?       ��  CDiodeBehavior     � ����        ��������� ���� 27     ��������� ����       ��������� ����       �������� D+D- j�     D+        ����D+����                        ��hd1n4007d1n4007               �hDiode   Generic   D1D1                D #�    ����D+D+      PASAA   ,����#�   ����D-D-      PASAK�d�����DiodeDiode	FairchildDO-41             10  j�    M-      ����M-����                        ��� 10  _10 	�    �    `   `   M+2  	�   j  `   �  M-3   �           IS1    	 �                    ��                                                               M+�                   ��                                                          �   M-�             <     ��     T                                                �     �       �     ��                                                        ̀ �����   @   <                  ����                                         ����<   @   �   � ����H   ����t     ��                                                        �  ������� �������  ��          @ @                                           �����x    ��b�����l    
>DA�����l    uT@ @ � ����D   <   |     ��                                                      ����D   <   |   ����D   <   |   [value]       �   �  �  Z     D   �   |   � ��������B        ��                                                       ��������B      ��������B      	[refname]       f   �    �     �����      
 ������  ���	   Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       Ԁ     � L	L�    �RS�-1.18m      �������� M+M- j�     M+        ����M+����                        ���AmmeterAmmeter   V            ��Analog Meters   Generic   IS1IS1          ����  VAm #�    ����M+M+      PASAM+�������#�   ����M-M-      PASAM-������Analog MetersAmmeter-verticalGeneric              3 �   |    �       _   �         _   �                 capacitor_generic�    x   �4 �	�    �       �   C-�  	�   �    �  �   C+�   �  �         C1     �                   ��                                                           @   C-�                   ��                                                      �   @   C+� �   @   `   @      ��    ��                                                � `   `   `         ��                                                        � @   `   @         ��    ��                                                � @   @       @     ��    p�H                                                �     `   �   �     ��                                                           `   �   �       `   �   �   [capacitance]       �     7  �      `   �   �   �         �   $     ��                                                               �   $           �   $   	[refname]       �  �  	  �          �   $    �����    �      ��   	Capacitor     Miscellaneous      �?       ��  CCapacitorBehavior     � '  -C��6?0.1m      ��������� ���� x     ��������� ����       ��������� ����       �������� C+C- j�     C+        ����C+����                        ��j�    C-      ����C-����                        �� 	capacitor   N           ��Passive   Generic   C1C1          ����  C #�    ����C+C+      PASAC+    ����#�   ����C-C-      PASAC-    ����Passive Generic              3  j�     M+        ����M+����                        ��[���  3   z 3 y 	�    �           M+i  	�   �   �     M-j   @              VRL    
 �                   ��                                                           `   M+�                   ��                                                      �   `   M-�     `       `     ��    ���                                                 � �   `   �   `     ��                                                       �    L      \     ��    ���                                                 �     T      T     ��    (�K                                                � �   X   �   X     ��               	FIXED_ROT                                        ̀     <   �   �                   ����                                             <   �   �   � (   D   �   x     ��                                                      (   D   �   x   (   D   �   x   [value]       �  �   �  Z  (   D   �   x   �        �   0    	 ��        	                                                      �   0          �   0   	[refname]       �  $   n  �          �   0    �  �����  ���      �
     	voltmeter    voltmeter_smallMiscellaneous      �?       ��   CVoltmeterBehavior     � ����   K,�-14.04      �������� M+M- �j�    M-      ����M-����                        ��	voltmeter	voltmeter   �            ��Analog Meters   Generic   VRLVRL          ����  IVm #�    ����M+M+      PASAM+- � ����#�   ����M-M-      PASAM-NAL
����Analog Meters Generic              4 � w ��  ��j�     M+        ����M+����                        ���  4   v 4 u 	�    �    `   `   M+2  	�   �   �
  �   �   ��   �
  @   � 	            	        `   �  M-3   �
           IS2    	 �                    ��                                                               M+�                   ��                                                          �   M-�             <     ��                                                        �     �       �     ��                                                        ̀ �����   @   <                  ����                                         ����<   @   �   � ����H   ����t     ��                                                        �  ������� �������  ��          @ @                                           �����x    ��b�����l    
>DA�����l    uT@ @ � ����D   <   |     ��                                                      ����D   <   |   ����D   <   |   [value]       T	  �  [
  Z     D   �   |   � ��������B        ��                                                       ��������B      ��������B      	[refname]       	  �  �	  �     �����      
 ������  ���	   Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       Ԁ     � ��9�    �BU�-1.30m      �������� M+M- �j�    M-      ����M-����                        ��AmmeterAmmeter   V            ��Analog Meters   Generic   IS2IS2          ����  VAm #�    ����M+M+      PASAM+LVIS����#�   ����M-M-      PASAM-TA
>����Analog MetersAmmeter-verticalGeneric              12 s  �j�     D+        ����D+����                        ��	 12  	 r 12 q 	�    �          D+   	�   �   �
  `	   �   ��   �
  �
   �                         @  D-    �
            D2     �                   ��                                                           `   D+�                   ��                                                          �   D-�     �       �      ��                                                        �     �   �����     ��                                                        �     �   �����     ��    .I @                                                �     `       �     ��    }͇0                                                �    �       �     ��    NDDA                                                �     �   �����     ��    G5                                                  �     �       �     ��     ��8                                                � 0   `   �   �    	 ��        	                                               0   `   �   �   0   `   �   �   	[devname]        �������������������������      � 0   �   �   �    
 ��        
                                               0   �   �   �   0   �   �   �   	[refname]       p  �  �  �	  ����   �   <    �������    ��          �� �  diode     Miscellaneous      �?       z�     � ����        ��������� ���� 27     ��������� ����       ��������� ����       �������� D+D- �j�    D-      ����D-����                        ��d1n4007d1n4007               ��Diode   Generic   D2D2                D #�    ����D+D+      PASAA�� ����#�   ����D-D-      PASAK � ����DiodeDiode	FairchildDO-41             11  j�     1       ����1����                        ��� 11   n 11 m �   L    n 0 �      n VControl 	�    �   �      1S  	�   \   �   �  2T  	�   ^       �  3U  	�             4V    
  `	       X4     �                    ��                                                       @   `   1�                   ��                                                      @   �   2�                   ��                                                          �   3�                   ��                                                          `   4�     �       `     ��    ��                                                �     �       �     ��                                                        �     �       �    
 ���   ��                                                � �����      �    	 ���   p�H                                                ��  TEllipse <   �   D   �                  ����                                         <   �   D   �   <   �   D   �   ̀ �����      �               	   ����                                         �����      �   � @   �   @   �     ��       
                                                � 0   �   @   �     ��    D�H                                                � @   �   @   `     ��                                                       �    �   �����     ��  � �H        	FIXED_ROT                                        �    �   4   �     ��    .I                                                  � `   �   �   �     ��                                                       `   �   �   �   `   �   �   �   	[refname]       @    �  �      (   t   L   � `   `   �   �     ��                                                       `   `   �   �   `   `   �   �   	[devname]        ����������������       �   (    ����      �  �	��     �  vcswitch     Miscellaneous      �?   9 
 >�    � ����      @4.5      ��������� ����      �?0.5     ��������� ����      �?0.5     ��������� ����    ��.A1meg     �������� 1234 �j�    2      ����2����                        ��j�    3      ����3����                        ��j�    4      ����4����                        ��X4_vcswitchX4_vcswitch
 9               �Switches   Generic   X4X4          ����B���voltage controlled switch   VCSW{.subckt vcsw 1 2 3 4
S 1 2 3 4 switch
.model switch sw (vt={(Von+Voff)/2} vh={(Von-Voff)/2} ron={Ron} roff={Roff})
.ends   D�    1turnon voltage   ParamSubVon               D�    1turnoff voltage   ParamSubVoffV             D�    0on resistance   ParamSubRonOhm             D�    0off resistance   ParamSubRoffOhm               X #�    ����11      PASA1H�~����#�   ����22      PASA2	   ����#�   ����33      PASA3�8  ����#�   ����44      PASA4�8  ����Switches Generic              0 ��   L    J 0 �    L     �           �   �           �   �               Gnd	�    �'   �  �   �   �   �  �                             `       Gnd}   `  �          gnd2     �                    ��                                                               Gnd�                   ��     �          AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��     5 (         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��    �׿         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         "#$&  %     Ground    
Ground DINMiscellaneous      �?       h�       Gnd j�     Gnd        ����Gnd����                        ��gndgnd                 (Analog Meters   Generic   gnd2gnd2          ����  gnd #�    ����GndGnd      GNDAGnd�����SourcesGroundGeneric              0 �   L     0  j�    V-      ����V-����                        ��k (+j�     1       ����1����                        ��j�    4      ����4����                        ��  0    J 0 fI 	�    T        �  1S  	�   n         2T  	�   *   �      3U  	�   b   �   �  4V   @  `	         X2     �                    ��                                                           �   1�                   ��                                                          `   2�                   ��                                                      @   `   3�                   ��                                                      @   �   4� @   �   @   �     ��    ��                                                � @   `   @   �     ��                                                        � @   �   @   �    
 ���   ��                                                � H   �   8   �    	 ���   p�H                                                 �    �   �����                  ����                                         �����      �   �����      �   ̀ P   �   0   �               	   ����                                         0   �   P   �   �     `       �     ��       
                                                �    �       �     ��    D�H                                                �     �       �     ��                                                       � 8   �   H   �     ��  � �H        	FIXED_ROT                                        � ,   �      �     ��                                                        � `   �   �   �     ��                                                       `   �   �   �   `   �   �   �   	[refname]       `    �  �  T   �   �   �   � �   �   @  �     ��                                                       `   `   �   �   `   `   �   �   	[devname]        ����������������T   `   �   �    2345;<>      7?  @9AB=68    : �  vcswitch     Miscellaneous      �?   9 
 >�    � ����      @4.5      ��������� ����      �?0.5     ��������� ����      �?0.5     ��������� ����    ��.A1meg     �������� 1234 ,gj�    3      ����3����                        ��-vcswitchvcswitch
 9               ,gH-Switches   Generic   X2X2          ����B���voltage controlled switch   VCSW{.subckt vcsw 1 2 3 4
S 1 2 3 4 switch
.model switch sw (vt={(Von+Voff)/2} vh={(Von-Voff)/2} ron={Ron} roff={Roff})
.ends   D�    1turnon voltage   ParamSubVon               D�    1turnoff voltage   ParamSubVoffV             D�    0on resistance   ParamSubRonOhm             D�    0off resistance   ParamSubRoffOhm               X #�    ����11      PASA1�S����#�   ����22      PASA2    ����#�   ����33      PASA3�U����#�   ����44      PASA4531E����Switches Generic              VControl � j�     V+        ����V+����                        ��" H5 G  VControl    VControl *	�    <           V+g  	�   !      �  V-h   �   	         VCtrl     �                   ��                                                           `   V+�                   ��                                                          �   V- �     �   �����                   ����                                         �����       �   �����       �   �    �   �����     ��    ��)                                                �     �       �     ��    ��`                                                �     �       �     ��    ��)                                                �     \       �     ��    p�Z                                                � �����   
   �    
 ��               	FIXED_ROT                                        � \   `   \   `     ��                                                      \   `   \   `   \   `   \   `           �   
  �   
                � 0   �   �   �     ��        	                                               0   �   �   �   0   �   �   �   [dc]       P  �
  ~  >          p   @   � 0   \   �   �    	 ��        
                                               0   \   �   �   0   \   �   �   	[refname]       P  
  @  �
      ����t       W  XY[VZ]^_      \    U �  Voltage Source    Voltage Source DINRoot      �?       ��  CVSourceBehavior     � ����        0      ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       �������� V+V- R+volt_sourcevolt_source   +0            R+Sources   Generic   VCtrlVCtrl          ����       �0����      $�-10      ���������0����      $@10     ���������0            0     ���������0��- a2U0*�3?300u     ���������0��- a2U0*�3?300u     ���������0@x}{�G�zd?2.5m     ���������0���{�G�zt?5m     ��������    �0            0      ���������0����      @5     ���������0����     �f@180     ���������0            0     ���������0            0     ��������    �0            0      ���������0����      �?1     ���������0����      �?1     ���������0            0     ���������0����      �?1     ��������    �0            0      ���������0����      �?1     ���������0            0     ���������0 N  �����>2u     ���������0'  ���ư>1u     ���������0'  ���ư>1u     ��������    �  ���� 0 0      ��������                0      �������� ����       �������� ����       �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������               V #�    ����V+V+      PWR+AV+NDDA����#�   ����V-V-      PWR-AV- � ����Sources Generic              z N  J & 8 � �� n _v cr � ~ �        L  � | x ep at � 0 ' 0                 � �  � � � ]    � �[ � � _ W �Y � ; � � � a U � Q � � � � � ) � � � � mS = 5 =     !T n��   � � � ^    � � � ��l` j��   \  < �   � � � � P � V X � � Z � � b � R � * ( : �   � � � � �      ��  CLetter    CEn el model real, els dos inductors estar�n acoplats magn�ticament.�  W    |      ����Arial����                       Arial     ��   �La tensi� de sortida puja una mica m�s si tenim diodes que converteixen el interruptors en interruptor unidireccionals, que no permeten que la corrent vagi cam a la font.�  �  J  �	      ����Arial����                       Arial     ��   oLa freq��ncia de traball ha d'estar molt ben ajustada a la freq. de resonancia de les bobines y el condensador.R  �  o  �      ����Arial����                       Arial     ��   ;Ajustant el temps en ON podem ajustar la tensi� de sortida.;  s  �        ����Arial����                       Arial     ��   dLa freq��ncia de treball ha de ser lleugerement superior a la corresponent a la freq. de resonancia.1  �  G  �      ����Arial����                       Arial     ��   �.Aquest dispositiu pot tenir un rendiment espant�s, tot i que se suposa un oscilador no a de tenir gaire consum.
Aix� sembla ser degut al desfase entre la tensi� de cuadrada y la filtrada.
Per solventar aquest desfase la conmutaci� ha d'estar sincronitzada amb la tensi� filtrada, no a un clock fix.
  �  �  z      ����Arial����                       Arial            
 �@ ����        ���������             0     ��������� ����      @5     ���������  ʚ;�������?.1     ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ���� true
     ��������� ����  false     ��������               
                  � ����        ��������� ����       ���������  ����       ���������@ ����       ���������@ ����       ��������               
                  � ����        ��������� ����       ���������@ ����       ���������  ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������               
                 � ����dec     ��������� ����     @�@1k     ��������� ����    ��.A1meg     ��������� ����       20     ��������� ���� true     ��������� ���� true     ��������� ���� true	     ��������� ����  false
     ��������               
                 �  ����        ���������  ����       ���������  ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����  	     ��������� ����  
     ��������               
                  	 � ����        ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������               
                 � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                    �             0      ���������  ʚ;�������?100m     ��������� �� �h㈵��>0.01m     ��������� �� �h㈵��>0.01m     ��������� ���� True     ��������� ����  F     ��������� ���� true     ��������� ����  false     ��������               
                 � ����     @�@1K      ���������  ����       ���������  ����       ���������  ����       ��������               
         ��              �  ����        ��������              
                  �  ����        ��������              
                                  
                 �@ ����        ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ���� true	     ��������� ����  false
     ��������� ���� true     ��������� ����  false     ��������               
                 � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                        � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                 � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                 � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                 �@ ����        ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����decade     ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������               
                 � ����        ��������� ����       ���������@ ����       ���������  ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������               
                        � ����dec     ��������� ����     @�@1k     ��������� ����    ��.A1meg     ��������� ����       20     ��������� ����        0     ��������� ����        0     ��������� ���� true	     ��������� ���� true
     ��������� ����      I@50     ��������� ���� true     ��������� ����  false     ��������               
                         / � ���� x'     ���������     �-���q=1E-12     ��������� @B -C��6?1E-4     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x	     ��������� ���� x!     ��������� ����    �  500
     ��������� ���� x     ��������� ����    �  500     ��������� ���� x$     ��������� ���� x$     ��������� ���� x%     ��������� ���� x"     ���������  ���� x*     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x&     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x+     ��������� ���� x,     ��������� ���� x-     ��������� ���� xg     ��������� ���� xf     ��������� ���� xd     ��������� ���� xe     ��������� ���� xh     ��������� ���� xj     ��������� ���� xi     ��������� ���� xk     ��������� ����    e��A1Gl     ���������             0�     ��������� ����      @5�     ��������� ����      @2.5�     ��������� ����      �?.5�     ��������� ����      @4.5�     ��������� 
   ��&�.>1n�     ��������� 
   ��&�.>1n�     ��������� 
   ��&�.>1n�     ��������� 
   ��&�.>1n�     ��������           ��  CPrimitiveModel    d1n4007   �    1�a��%>2.55e-9      ��������� ���� 27     ���������  �/�$��?0.042     ��������� ����      �?1.75     ���������  �  ��v��(�>5.76e-6     ���������     �]}IW�=1.85e-11     ��������� ����      �?0.75     ��������� ����Zd;�O�?0.333     ��������� ���� 1.11	     ��������� ���� 3.0
     ���������      0     ��������� ���� 1     ��������� ���� 0.5     ��������� ����     @�@1000     ��������� � Ǯ���?9.86e-5     ��������     Diode Generic��   CPrimitiveModelType Junction Diode model����DD   D����� 1.0E-14Saturation current    ProcessisAmp0       e     D����� 27!Parameter measurement temperature    ProcesstnomDeg C0     s     D����� 0Ohmic resistance    ProcessrsOhm0      f     D����� 1Emission Coefficient    Processn 0      g     D����� 0Transit Time    Processttsec0     h     D����� 0Junction capacitance    ProcesscjoF0     i     D����� 0     Processcj0F0     i     D����� 1Junction potential    ProcessvjV0      j     D����� 0.5Grading coefficient    Processm 0      k     D����� 1.11Activation energy    ProcessegeV0     	 l     D����� 3.0#Saturation current temperature exp.    Processxti 0     
 m     D����� 0flicker noise coefficient    Processkf 0      t     D����� 1flicker noise exponent    Processaf 0      u     D����� 0.5#Forward bias junction fit parameter    Processfc 0      n     D����� infReverse breakdown voltage    ProcessbvV0      o     D����� 1.0e-3$Current at reverse breakdown voltage    ProcessibvA0      p     D�����  Ohmic conductance    ProcesscondMho     r        D��     ?C
                Ariald     h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j                   ����            (�T               ��  TSignal                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                      v(vrl)       ����                  ȃ                     
i(isource)       ����                  ȃ                     i(is1)       ����                  ȃ                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CDCsweep       
 ����������               
                       ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                       v(vrl)       ����                  ȃ                      
i(isource)       ����                  ȃ                      i(is1)       ����                  ȃ                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACsweep        ��������               
                       ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                      v(vrl)       ����                  ȃ                     
i(isource)       ����                  ȃ                     i(is1)       ����                  ȃ                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  �� 
 CTranSweep       ��������               
                       ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                       v(vrl)       ����                  ȃ                      
i(isource)       ����                  ȃ                      i(is1)       ����                  ȃ                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACdisto        �����               
                           ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                       v(vrl)       ����                  ȃ                      
i(isource)       ����                  ȃ                      i(is1)       ����                  ȃ                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  �        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                           ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                       v(vrl)       ����                  ȃ                      
i(isource)       ����                  ȃ                      i(is1)       ����                  ȃ                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  �        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                           ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                       v(vrl)       ����                  ȃ                      
i(isource)       ����                  ȃ                      i(is1)       ����                  ȃ                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  �        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                           ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                       v(vrl)       ����                  ȃ                      
i(isource)       ����                  ȃ                      i(is1)       ����                  ȃ                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  �        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                           ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                       v(vrl)       ����                  ȃ                      
i(isource)       ����                  ȃ                      i(is1)       ����                  ȃ                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  �        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
         �             	    ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                      v(vrl)       ����                  ȃ                     
i(isource)       ����                  ȃ                     i(is1)       ����                  ȃ                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACnoise        ��������               
                    
    ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                      v(vrl)       ����                  ȃ                     
i(isource)       ����                  ȃ                     i(is1)       ����                  ȃ                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��         �  ����        ���������  ����       ���������  ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����  	     ��������� ����  
     ��������              
                        ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                      v(vrl)       ����                  ȃ                     
i(isource)       ����                  ȃ                     i(is1)       ����                  ȃ                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CFourier        ����               
         ��                   ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                      v(vrl)       ����                  ȃ                     
i(isource)       ����                  ȃ                     i(is1)       ����                  ȃ                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACpz        	 ���������               
                       ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                      v(vrl)       ����                  ȃ                     
i(isource)       ����                  ȃ                     i(is1)       ����                  ȃ                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CDCtf         �����               
                       ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                      v(vrl)       ����                  ȃ                     
i(isource)       ����                  ȃ                     i(is1)       ����                  ȃ                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CDCsens         �����������               
                       ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                       v(vrl)       ����                  ȃ                      
i(isource)       ����                  ȃ                      i(is1)       ����                  ȃ                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j                  ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                      v(vrl)       ����                  ȃ                     
i(isource)       ����                  ȃ                     i(is1)       ����                  ȃ                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CShow         �              
                       ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                      v(vrl)       ����                  ȃ                     
i(isource)       ����                  ȃ                     i(is1)       ����                  ȃ                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CShowmod         �              
                       ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                      v(vrl)       ����                  ȃ                     
i(isource)       ����                  ȃ                     i(is1)       ����                  ȃ                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  �� 
 CLinearize        �  ����        ��������               
                       ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                      v(vrl)       ����                  ȃ                     
i(isource)       ����                  ȃ                     i(is1)       ����                  ȃ                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CParamTranSweep        �������������               
                       ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                      v(vrl)       ����                  ȃ                     
i(isource)       ����                  ȃ                     i(is1)       ����                  ȃ                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  �              ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                       v(vrl)       ����                  ȃ                      
i(isource)       ����                  ȃ                      i(is1)       ����                  ȃ                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CParamACSweep        RSTUVWXYZ[\]^               
                       ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                      v(vrl)       ����                  ȃ                     
i(isource)       ����                  ȃ                     i(is1)       ����                  ȃ                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CMonteCarlo_op        ����������������������������               
                              ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                      v(vrl)       ����                  ȃ                     
i(isource)       ����                  ȃ                     i(is1)       ����                  ȃ                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CMonteCarlo_dc        �� 	
               
                       ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                       v(vrl)       ����                  ȃ                      
i(isource)       ����                  ȃ                      i(is1)       ����                  ȃ                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CMonteCarlo_ac         !"#$%&'()*+,-./012345               
                       ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                      v(vrl)       ����                  ȃ                     
i(isource)       ����                  ȃ                     i(is1)       ����                  ȃ                     i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CMonteCarlo_tran        6789:;<=>?@ABCDEFGHIJKLMNOPQ               
                       ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                       v(vrl)       ����                  ȃ                      
i(isource)       ����                  ȃ                      i(is1)       ����                  ȃ                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CACsens        _`abcdefghi               
                              ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                       v(vrl)       ����                  ȃ                      
i(isource)       ����                  ȃ                      i(is1)       ����                  ȃ                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j  ��  CNetworkAnalysis        jklmnopqrst               
                       ����            P               ȃ                        v(vcontrol)       ����                  ȃ                       
v(vsource)       ����                  ȃ                       v(3)       ����                  ȃ                       v(4)       ����                  ȃ                       v(6)       ����                  ȃ                       v(7)       ����                  ȃ                       v(11)       ����                  ȃ                       v(10)       ����                  ȃ                       v(12)       ����                  ȃ	                       v(13)       ����                  ȃ
                       i(vctrl)       ����                  ȃ                       v(vrl)       ����                  ȃ                      
i(isource)       ����                  ȃ                      i(is1)       ����                  ȃ                      i(is2)       ����                  h�  �� �|p�|����m�|+j  h�  �� �|p�|����m�|+j                  ����            P              33�=           ��   CDigSimResTemplate                ���       ����  ����:�0�yU>20.00n���   ����                       Arial����                       Arial����                       Arial  �   �  �                                ����  ���� ������       ����  ���� ������                 �               ����  �����       200������         0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial      �       �         �     �   �  �  Circuit1                  ����  ��    ��������                                                                                                                                                                                                                                 g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     ��   CPackageAliasSuperPCBStandardDIODE3      ΅Eagle	DIODE.LBRDO41-7   AC  ΅Orcad 	DAX2/DO41      ΅	Ultiboard	L7DIO.l55DIO_DO41              A      g   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     ����        A                                            �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            J  �                L L�� �� C KE                 2         �  �              � � �           ����    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                      �  �                ̀         �  @                  ���                                                  �  @  �     <   �  <     ��                                                        �     |   �  |     ��                                                        �     �   �  �     ��                                                        �     �   �  �     ��                                                        � �      �  4     ��                                                      �      �  4   �      �  4   [title]                                       � �   D   �  t     ��                                                      �   D   �  t   �   D   �  t   [description]                                       � `   �   h  �     ��                                                      `   �   h  �   `   �   h  �   [id]                                       � �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       �      �   8    ��        	                                                   �   8       �   8  Date :       �    8
  �                  � �     �  4   	 ��        
                                              �     �  4  �     �  4  [date]                                       �       t   8    
 ��                                                            t   8         t   8   Title :       �    
  �                  �    L   �   x     ��                                                         L   �   x      L   �   x   Description :       �  �  �  �                  �    �   �   �     ��                                                         �   �   �      �   �   �   ID :       �  �  �	  T                  �    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �  L  (                     ��������������          �     	title box    Analog Misc      �?    9 
 >�     �  ����        ���������  ����       ���������  ����       ���������  ����       ���������  ����       ��������        9                                      ����B��� ����     D�            title                D�            description               D�            id               D�            designer               D�            date                           ����            `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                                                                                            2         �  �              � � �                   ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                          �   ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    
cgs 76         47 80moh5.6  m = 0.3mvrd nmodel 00   ibv2.     ȃ                      TIME� # ) time                      ȃ                        v(3)      v(3)    TIME                 ȃ                        i(vctrl)� �   i(vctrl)    TIME                 ȃ                       v(vcontrol)      v(vcontrol)    TIME                 ȃ    (v(3)-v(4))                   v(VRL)� �   v(VRL)    TIME                 ȃ                       i(irl)�   � i(irl)    TIME                 ȃ                        v(4)      v(4)    TIME                 ȃ    i(irl)*v(vrl)                    PRL  � �  ����TIME                 ȃ                        
v(vsource)      
v(vsource)    TIME                 ȃ                       
i(isource)�   � 
i(isource)    TIME                 ȃ                      i(is1)  � � i(is1)    TIME                 ȃ                      i(is2)� �   i(is2)    TIME                 ȃ    i(isource)*v(vsource)                    PSource@ � �  ����TIME                 ȃ                        v(11)      v(11)    TIME                           2         �  �           Time  � � �               0     ����                       Arial����                       Arial                              ����  ������)��?6.915528e-002���A8)      ����  ������)��?6.915528e-002���A8)      ����  �����@M�?2.547151e-001������      ����  �����@M�?2.547151e-001������                                                                           �                      �                                                                                                                                                                                                                                                                  �  �                                                                                                                                                                                                                                                                              �  �                                                                                                                                                                                                                                                                                                                                                                  1m  0                            100   100                                                             1m  0                            100   100                                1m  0                            100   100                                1m  0                            100   100                                                 
                 1m  0                            100   100                            ��   CPartPackage     ��   CPackageg   DO-41�3 pin diode package                                                                                                                                                                                                                                       �     ����    �           ��   CMiniPartPin    ����V+V+     PWR+V+g      �   ����V-V-     PWR-V-h     voltage_sourcevoltage_source                          �    ����M+M+     PASM+i      �   ����M-M-     PASM-j     	voltmeter	voltmeter                          �    ����11     PAS1�      �   ����22     PAS2�     BatteryBattery                          �    ����GndGnd     GNDGnd}      GndGnd                  �    ����MM       ��������MarkerMarker                  �    ����GndGnd     GNDGnd}      GndGnd                  �    ����M+M+     PASM+2      �   ����M-M-     PASM-3     Ammeter2Ammeter2                          �    ����11     PAS1S      �   ����22     PAS2T     �   ����33     PAS3U     �   ����44     PAS4V     vcswitchvcswitch                                          �    ����MM       ��������MarkerMarker                  �    ����MM       ��������MarkerMarker                  �    ����L+L+     PASL+K      �   ����L-L-     PASL-L     InductorInductor                          �    ����C+C+     PASC+�      �   ����C-C-     PASC-�     capacitor_genericcapacitor_generic                          �    ����L+L+     PASL+K      �   ����L-L-     PASL-L     InductorInductor                          �    ����11     PAS1S      �   ����22     PAS2T     �   ����33     PAS3U     �   ����44     PAS4V     vcswitchvcswitch                                          �    ����M+M+     PASM+2      �   ����M-M-     PASM-3     Ammeter2Ammeter2                          �    ����M+M+     PASM+2      �   ����M-M-     PASM-3     Ammeter2Ammeter2                        �    ����D+D+     PASA       �   ����D-D-     PASK       c  ��   CPackagePin 1 D+PAS  AA'� 2 D-PAS  AKDiodeDiode	Fairchild      1n4007 D1n4007D1            diode-21n40071n4007                        �    ����D+D+     PASA       �   ����D-D-     PASK       r   '� 1 D+PAS  AA'� 2 D-PAS  AKDiodeDiode	Fairchild      1n4007 D1n4007D2            diode-21n40071n4007                          �    ����R+R+     PASR+  �,  �   ����R-R-     PASR-  �,  resistor_genericresistor_generic                          �    ����M+M+     PASM+0  �  �   ����M-M-     PASM-1  �  AmmeterAmmeter                          �    ����MM       ��������MarkerMarker                                                                                                                                                                                                                                                                                                    
m1     8 8 mm l=100u w                        used                             ��    �����Z��� ��                        X�T                                                                                                                                                           `                               �i��    �i��     � ����                        ���                                   �&��0�u .I �   �                         �                                                                                                                                                                                       ���    �����������                            �i��                            ��               �����                        �@�                            �i��    �i�������@
KCTRL                        ���                            ?Q    �?Q�?Q@QXP                        �P                            Ha    �_\PU�_\`\                        c\                            TRL.      
QVI_SOURCE.I                         G5                              �[�    h\��\��\�0]�                        `�X                            ×sA    S1.I Le�7
JL2.I                         G6                                                                                                         
G5    A
G4 =���
G3 5�                        A
>D                            �T    (T��U�U �U                        �V                                                                                                            �C�?    �W�dV �  �                          ��    2 2 2 2 d                                                                                 