    � B2SPICE zzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz    ��  CPart    �����   �  �  �����   �  �              voltage_source��  CIntPin    ��  CWire    �        �
   /   �   �      /   �   �                  Marker ��  CExtPin    ��  CVertex
   �  `   ��  CSegment    �   �  �                    
        `      M     @  @          Ctrl1     ��   CPin                   ��                                                           `   M��  TLine     P       `     ��    ��                                                ��  TPolygon     ����    ����   ��                                                         ��  TPoint    0        �   @        �    P        �0   @            ��  
 TTextField    �����        ��                                                          �����         �����      	[refname]       X  1  0  �        �   ,               Marker     Miscellaneous      �?    +   ��   CMarkerBehavior     ��  CValue             0.0      �������� M ��  	 TModelPin ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �         �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               " Analog MiscV   Generic   Ctrl1Ctrl1          ����               Ctrl1  v(Ctrl1)  N ��   CPartPin    ����MM       A     ����RootmarkerGeneric              Ctrl1 �        �   /   �   �      /   �   �                  Marker% 	�    �    @  �   �   ( �   @  �   )                       `      MȘ� �
  `          Ctrl1     �                   ��                                                           `   M�     P       `     ��                                                        �     ����    ����   ��                                                         �    0        �   @        �    P        �0   @            �    �����        ��                                                          �����         �����      	[refname]       �
  Q  �  �        �   ,    -   + 2 ,      Marker     Miscellaneous      �?    +   �     �             0.0      �������� M !� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      3   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               5 Analog MiscV   Generic   Ctrl1Ctrl1          ����               Ctrl1  v(Ctrl1)  N #�    ����MM       A  �����RootmarkerGeneric              Ctrl1 �        �   /   �   �      /   �   �                  Marker7 	�    �       	   �   : �      `	   ;                       `      M���� �  �          Ctrl1     �                   ��                                                           `   M�     P       `     ��     �                                                 �     ����    ����   ��                                                         �    0        �   @        �    P        �0   @            �    �����        ��                                                          �����         �����      	[refname]       �  �  �  q        �   ,    ?   = D >      Marker     Miscellaneous      �?    +   �     �             0.0      �������� M !� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �      E   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               G Analog MiscV   Generic   Ctrl1Ctrl1          ����               Ctrl1  v(Ctrl1)  N #�    ����MM       A �������RootmarkerGeneric              Ctrl1 �      �       �   �  �      �   �  �              vcswitch�    �     �    L     �           �   �           �   �               GndM 	�    �   �      �   �   �      �   �   �  �
   S         R     Q      P     �   P �   �
      �   �*   �
  �
   W          V     U          �   �   �  �
   Y          P                 `       Gnd}   `             gnd1     �                    ��                                                               Gnd�                   ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��    ��)         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��    p�Z         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         [ \ ] _   ^      Ground    
Ground DINMiscellaneous      �?       ��   CGroundBehavior       Gnd ��   CBehPin     Gnd        ����Gnd����                        ��gndgnd                 c Analog Meters   Generic   gnd1gnd1          ����  gnd #�    ����GndGnd      GNDAGnd �)����SourcesGroundGeneric              0 �   L    �           �   �          �   �              Battery�    �    g �    h    �       _   @  �      _   @  �              Ammeter2i �   �    �   l   �       �   �  �      �   �  �              vcswitch�    �    o �   p   �       �   �  �      �   �  �              	voltmeter�    �    �   t   �       �   �  �       �   �  �               R�    p    v 3 u 	�    �   `	  �   �
   y �   �
  �   z �   �   �
      �   �    
      ~        }     �   �   �
  `   �         }     |     {     �   { �)   �
  `	   �                               �  �   R+  	�   �   �  �   �	   �	   �  �   � �   �   �      �   � �   �      �             �   �$   �  `   �         �     �     �     �   � �   �  `	   �                �                  �   R-   �  �         R     �                    ��                                                       �   @   R+�                   ��                                                          @   R-�    @   $   0     ��    ��)                                                � 0   P   $   0     ��                                                        � 0   P   <   0     ��    ��)                                                � H   P   <   0     ��    p�Z                                                � H   P   T   0     ��                                                       � `   P   h   @     ��    D�Z                                                � �   @   h   @     ��    ��d                                                � `   P   T   0    	 ��    |�f	                                                �    @       @    
 ��    <�b
                                                �     `   �   �     ��                                                           `   �   �       `   �   �   [resistance]       �   	  P  �	      `   �   �   �         t   $     ��                                                               t   $           t   $   	[refname]       �  �  (  �          t   $    � � � � � � � � � � � � �    resistor    resistor DINMiscellaneous      �?       ��  CResistorBehavior     � ����      6@22      ��������� ���� 27     ��������� ����       ��������� ����       �������� R+R- b�     R+        ����R+����                        ��b�    R-      ����R-����                        �� resistor                � � Passive   Generic   RR          ����    R #�    ����R+R+      PASAR+JV1.����#�   ����R-R-      PASAR-�)����Passivedefault resistor, 1KGeneric              6 s �    t    �       �   �  �      �   �  �              vcswitch� �   l   � 5 �   �    �    �    �   /   �   �      /   �   �                  Marker� 	�    �&      �   �   � �"      �   �                       `      M� �  `          Ctrl2     �                   ��                                                           `   M�     P       `     ��     �                                                 �     ����    ����   ��                                                         �    0        �   @        �    P        �0   @            �    �����        ��                                                          �����         �����      	[refname]       �  Q  �  �        �   ,    �   � � �      Marker     Miscellaneous      �?    +   �     �             0.0      �������� M !� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               � Analog MiscV   Generic   Ctrl2Ctrl2          ����               Ctrl2  v(Ctrl2)  N #�    ����MM       A zzzz����RootmarkerGeneric              Ctrl2 �    �    �   /   �   �      /   �   �                  Marker� 	�    �   @   	   �   � �!   @  `	   �                       `      Mhz� �
  �          Ctrl2     �                   ��                                                           `   M�     P       `     ��                                                        �     ����    ����   ��                                                         �    0        �   @        �    P        �0   @            �    �����        ��                                                          �����         �����      	[refname]       �
  �  �  q        �   ,    �   � � �      Marker     Miscellaneous      �?    +   �     �             0.0      �������� M !� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               � Analog MiscV   Generic   Ctrl2Ctrl2          ����               Ctrl2  v(Ctrl2)  N #�    ����MM       A pH�����RootmarkerGeneric              Ctrl2 �    �    �   /   �   �      /   �   �                  Marker� 	�    �%   �  `   �    � �+   �  �   �                        `      MG5   �  @          Ctrl2     �                   ��                                                           `   M�     P       `     ��    �@
                                                �     ����    ����   ��                                                         �    0        �   @        �    P        �0   @            �    �����        ��                                                          �����         �����      	[refname]       �  1  p  �        �   ,    �   � � �      Marker     Miscellaneous      �?    +   �     �             0.0      �������� M !� ����M����        M����                                         0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    ��������             0��    �������� d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������                             ����  ����:�0�yE>10e-9��d         ����  ����:�0�yE>10e-9��d   �     � �   �����     ��   d   :�0�yE>10e-9��    �������� d   :�0�yE>10e-9��    ��������MarkerMarker  +               � Analog MiscV   Generic   Ctrl2Ctrl2          ����               Ctrl2  v(Ctrl2)  N #�    ����MM       A �����RootmarkerGeneric              Ctrl2 �    �    �   �����   �  �  �����   �  �              voltage_source� �   L    � 0 	�    �           V+g  	�   �'   �  @   �   � �   �  �   �                            �  V-h   �  �         V2     �                   ��                                                           `   V+�                   ��                                                          �   V-��  TEllipse     �   �����                   ����                                         �����       �   �����       �   �    �   �����     ��                                                        �     �       �     ��    1.I                                                 �     �       �     ��    G4                                                  �     \       �     ��    .I                                                 � �����   
   �    
 ��    G3 �        	FIXED_ROT                                        � \   `   \   `     ��                                                      \   `   \   `   \   `   \   `           �  �  �  �                � 0   �   �   �     ��        	                                               0   �   �   �   0   �   �   �   [dc]       p  P  �  �          p   @   � 0   \   �   �    	 ��        
                                               0   \   �   �   0   \   �   �   	[refname]       p  �  �  T      ����t       �   � � � � � � � �       �     �  �  Voltage Source    Voltage Source DINRoot      �?       ��  CVSourceBehavior     � ����        0      ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       �������� V+V- b�     V+        ����V+����                        ��b�    V-      ����V-����                        ��volt_sourcevolt_source   +0            Sources   Generic   V2V2          ����       �0����      @5      ���������0            0     ���������0            0     ���������0��� ����MbP?1m     ���������0��� ����MbP?1m     ���������0���{�G�zt?5m     ���������0 '�~j�t��?12m     ��������    �0            0      ���������0����      @5     ���������0����     ��@10k     ���������0            0     ���������0            0     ��������    �0            0      ���������0����      �?1     ���������0����      �?1     ���������0            0     ���������0����      �?1     ��������    �0            0      ���������0����      �?1     ���������0            0     ���������0 N  �����>2u     ���������0'  ���ư>1u     ���������0'  ���ư>1u     ��������    �  ���� 0 0      ��������                0      �������� ����       �������� ����       �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������               V #�    ����V+V+      PWR+AV+ �@
����#�   ����V-V-      PWR-AV-    ����Sources Generic              Ctrl2 �   �   �       �   �  �      �   �  �              vcswitch�    L     !0 �   p   !3  �   L    !0 	�    X        �  1S  	�   �          2T  	�   �   �      3U  	�   �   @  �
                   �   �  4V   �
  @         X6     �                    ��                                                           �   1�                   ��                                                          `   2�                   ��                                                      @   `   3�                   ��                                                      @   �   4� @   �   @   �     ��    ��                                                � @   `   @   �     ��                                                        � @   �   @   �    
 ���   ��                                                � H   �   8   �    	 ���   p�H                                                �    �   �����                  ����                                         �����      �   �����      �   �� 
 TRectangle P   �   0   �               	   ����                                         0   �   P   �   �     `       �     ��       
                                                �    �       �     ��    D�H                                                �     �       �     ��                                                       � 8   �   H   �     ��  � �H        	FIXED_ROT                                        � ,   �      �     ��                                                        � `   �   �   �     ��                                                       `   �   �   �   `   �   �   �   	[refname]       �  �	    �
      (   t   L   � `   `   �   �     ��                                                       `   `   �   �   `   `   �   �   	[devname]        ����������������       �   (    *+,-457      /8  91:;6.0    2 �  vcswitch     Miscellaneous      �?   9 
 ��  CParamSubBehavior    � ����������@4.9      ��������� �����������?1.1     ��������� ����      �?0.5     ��������� ����    ��.A1meg     �������� 1234 b�     1       ����1����                        ��b�    2      ����2����                        ��b�    3      ����3����                        ��b�    4      ����4����                        ��X6_vcswitchX6_vcswitch
 9               BCDESwitches   Generic   X4X4          ������   CParamSubModelType��voltage controlled switch   VCSW{.subckt vcsw 1 2 3 4
S 1 2 3 4 switch
.model switch sw (vt={(Von+Voff)/2} vh={(Von-Voff)/2} ron={Ron} roff={Roff})
.ends   ��  	 CParmDefn    1turnon voltage   ParamSubVon               H�    1turnoff voltage   ParamSubVoffV             H�    0on resistance   ParamSubRonOhm             H�    0off resistance   ParamSubRoffOhm               X #�    ����11      PASA1O�����#�   ����22      PASA2    ����#�   ����33      PASA3    ����#�   ����44      PASA4�XQ����Switches Generic              Ctrl2 �  � D� �  Ctrl2  � Ctrl2 �   L    � 0 	�    �    �   �  1S  	�   �#   �  �   �   �-   �  @   �   �,   �
  @   W�   X�   �
  �   Y               V    �   �(   �  @   �   \�   �  �   ]           [    V    U    T             �      2T  	�   �          3U  	�   �      `                       �  4V      �        X4     �                    ��                                                       @   �   1�                   ��                                                      @   `   2�                   ��                                                          `   3�                   ��                                                          �   4�     �       �     ��                                                        �     `       �     ��                                                        �     �       �    
 ���                                                       � �����      �    	 ���                                                       � D   �   <   �                  ����                                         <   �   D   �   <   �   D   �   3�    �   �����               	   ����                                         �����      �   � @   `   @   �     ��        
                                                � 0   �   @   �     ��                                                        � @   �   @   �     ��                                                        �    �   �����     ��  �             	FIXED_ROT                                        �    �   4   �     ��                                                        � `   �   �   �     ��                                                       `   �   �   �   `   �   �   �   	[refname]          |  �        (   t   L   �     �  <    ��                                                       `   `   �   �   `   `   �   �   	[devname]        ����������������       �   (    bcdekln      go  piqrmfh    j �  vcswitch     Miscellaneous      �?   9 
 =  X #�    ����11      PASA1G1  ����#�   ����22      PASA2VA_I����#�   ����33      PASA3�2�����#�   ����44      PASA4d   ����Switches Generic              6 �   t   J 6  � b�     M+        ����M+����                        ��b�    2      ����2����                        ��B 6   r 6 q 	�    �           M+i  	�      �     M-j   �             IV_VRL    
 �                   ��                                                           `   M+�                   ��                                                      �   `   M-�     `       `     ��    ��                                                � �   `   �   `     ��                                                        �    L      \     ��    ��                                                �     T      T     ��    p�H                                                � �   X   �   X     ��               	FIXED_ROT                                        3�     <   �   �                   ����                                             <   �   �   � (   D   �   x     ��                                                      (   D   �   x   (   D   �   x   [value]       �  �  �  b  (   D   �   x   �        �   0    	 ��        	                                                      �   0          �   0   	[refname]       �  $  @	  �         �   0    �  |}~��  ���      
     	voltmeter    voltmeter_smallMiscellaneous      �?       ��   CVoltmeterBehavior     � ����  ��b!@ 4.78      �������� M+M- xb�    M-      ����M-����                        ��	voltmeter	voltmeter   _            x�Analog Meters   Generic   IV_VRLIV_VRL          ����  IVm #�    ����M+M+      PASAM+    ����#�   ����M-M-      PASAM-    ����Analog Meters Generic              3 w # b�     1       ����1����                        ��� �C 3   n 3 m �      n Ctrl1 �   L    n 0 	�    �        �  1S  	�   Z         2T  	�   *   �      3U  	�   �    @  `                   �   �  4V   �
  �         X3     �                    ��                                                           �   1�                   ��                                                          `   2�                   ��                                                      @   `   3�                   ��                                                      @   �   4� @   �   @   �     ��                                                        � @   `   @   �     ��                                                        � @   �   @   �    
 ���                                                       � H   �   8   �    	 ���                                                       �    �   �����                  ����                                         �����      �   �����      �   3� P   �   0   �               	   ����                                         0   �   P   �   �     `       �     ��    D�H
                                                �    �       �     ��                                                       �     �       �     ��                                                        � 8   �   H   �     ��  �             	FIXED_ROT                                        � ,   �      �     ��                                                        � `   �   �   �     ��                                                       `   �   �   �   `   �   �   �   	[refname]       �  |          (   t   L   �     �  <    ��                                                       `   `   �   �   `   `   �   �   	[devname]        ����������������       �   (    �������      ��  �������    � �  vcswitch     Miscellaneous      �?   9 
 <�    � ����������@4.9      ��������� �����������?1.1     ��������� ����      �?0.5     ��������� ����    ��.A1meg     �������� 1234 �yb�    3      ����3����                        ��b�    4      ����4����                        ��vcswitchvcswitch
 9               �y��Switches   Generic   X3X3          ����F���voltage controlled switch   VCSW{.subckt vcsw 1 2 3 4
S 1 2 3 4 switch
.model switch sw (vt={(Von+Voff)/2} vh={(Von-Voff)/2} ron={Ron} roff={Roff})
.ends   H�    1turnon voltage   ParamSubVon               H�    1turnoff voltage   ParamSubVoffV             H�    0on resistance   ParamSubRonOhm             H�    0off resistance   ParamSubRoffOhm               X #�    ����11      PASA1  �����#�   ����22      PASA2  � ����#�   ����33      PASA3    ����#�   ����44      PASA4    ����Switches Generic              5 k �  yb�    M-      ����M-����                        ��C 5  j 5 	�    �   �   	   �   ��   �  `	   �                       `   �  M+2  	�   ^  `   `   M-3   @            VA_Ix1    	 �                    ��                                                           �   M+�                   ��                                                              M-�     �       �     ��                                                        �     <             ��                                                        3� @   <   �����                  ����                                         ����<   @   �   � ����x   ����L     ��                                                        �  ������� �������  ��          @ @                                           �����H    ��b�����T    
>DA�����T    uT@ @ � ����D   <   |     ��                                                      ����D   <   |   ����D   <   |   [value]         �  �  �     D   �   |   � ��������O        ��                                                       ��������O      ��������O      	[refname]       �   �  =  �     �����      
 ������  ���	   Ammeter-Vert    Ammeter-vert_smallMiscellaneous      �?       ��   CAmmeterBehavior     � ����   ����?217.40m      �������� M+M- b�     M+        ����M+����                        ���AmmeterAmmeter   V            ��Analog Meters   Generic   VA_Ix1VA_Ix1          ����  VAm #�    ����M+M+      PASAM+��W����#�   ����M-M-      PASAM-8�W����Analog MetersAmmeter-verticalGeneric              4  b�     1       ����1����                        ��� 4   f 4 e 	�    �   `       1�  	�   T   `   �  2�   @  `	          X1     �                    ��                                                               1�                   ��                                                          �   2�             $     ��    ��)                                                �     \       �     ��                                                        �    8   0   8    	 ��    ��)                                                �     H   @   H     ��    p�Z                                                �     $   @   $     ��                                                       �    \   0   \     ��    D�Z                                                �               ���                                                      �               ���   �Z	                                                � `          $    
 ��        
                                               `          $   `          $   	[devname]        ����������������`          $   � `   $      H     ��                                                       `   $      H   `   $      H   	[refname]       `  �	  �  l
  `   $      H    ��������    ��    �  �     Battery     Miscellaneous      �?    9 
 <�     � ����      @5      �������� 12 �b�    2      ����2����                        ��BatteryBattery
 9 i             ��Sources   Generic   X1X1          ����F���    BATTERY2.SUBCKT Xbattery 1 2
V1 1 2 DC {voltage}
.ENDS
   H�    1battery voltage   ParamSubvoltageV                X #�    ����11      PASA1�1b����#�   ����22      PASA20Ab����SourcesBatteryGeneric              0 "K �    L     �           �   �           �   �               Gnd�	�    �   `       Gnd}   �
  `          gnd2     �                    ��                                                               Gnd�                   ��    ��         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         ����  �     Ground    
Ground DINMiscellaneous      �?       `�       Gnd b�     Gnd        ����Gnd����                        ��gndgnd                 �Analog Meters   Generic   gnd2gnd2          ����  gnd #�    ����GndGnd      GNDAGnd    ����SourcesGroundGeneric              0 ��    L     �	           �   �           �   �               Gnd�	�    �      �
            	        `       Gnd}   �  �
          gnd3     �                    ��                                                               Gnd�                   ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         ����  �     Ground    
Ground DINMiscellaneous      �?       `�       Gnd b�     Gnd        ����Gnd����                        ��gndgnd                 �Analog Meters   Generic   gnd3gnd3          ����  gnd #�    ����GndGnd      GNDAGnd    ����SourcesGroundGeneric              0 �   L    J 0 �    L     �           �   �           �   �               Gnd�	�    �   �  �   �   �   �  @   �         �                `       Gnd}   @  �          gnd4     �                    ��                                                               Gnd�                   ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��    D�H         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��    x�W         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��    X��         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ                Ground    
Ground DINMiscellaneous      �?       `�       Gnd b�     Gnd        ����Gnd����                        ��gndgnd                 Analog Meters   Generic   gnd4gnd4          ����  gnd #�    ����GndGnd      GNDAGnd    ����SourcesGroundGeneric              0 �   L     0 �    L     �           �   �           �   �               Gnd
	�    a   `       Gnd}   �  `          gnd5     �                    ��                                                               Gnd�                   ��    p�H         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��    D�H         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ                Ground    
Ground DINMiscellaneous      �?       `�       Gnd b�     Gnd        ����Gnd����                        ��gndgnd                 Analog Meters   Generic   gnd5gnd5          ����  gnd #�    ����GndGnd      GNDAGnd�����SourcesGroundGeneric              0 Q�    L     �           �   �           �   �               Gnd	�    )   `       Gnd}   �
  �
          gnd6     �                    ��                                                               Gnd�                   ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��       0         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��       �         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ                Ground    
Ground DINMiscellaneous      �?       `�       Gnd b�     Gnd        ����Gnd����                        ��gndgnd                 Analog Meters   Generic   gnd6gnd6          ����  gnd #�    ����GndGnd      GNDAGnd��������SourcesGroundGeneric              0 $�    L     �           �   �           �   �               Gnd 	�    �    `       Gnd}   �  �          gnd7     �                    ��                                                               Gnd�                   ��    �@
         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �         @         ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    ,   4   ,     ��                 AMJ     AMJ AMJ AMJ AMJ AMJ AMJ        �    8   (   8     ��    KCTR         AMJ     AMJ AMJ AMJ AMJ AMJ AMJ         #$%'  &     Ground    
Ground DINMiscellaneous      �?       `�       Gnd b�     Gnd        ����Gnd����                        ��gndgnd                 )Analog Meters   Generic   gnd7gnd7          ����  gnd #�    ����GndGnd      GNDAGnd    ����SourcesGroundGeneric              0 �  b�    V-      ����V-����                        ����c ���EB)  0    J 0 wI �	�    Z    �   �  1S  	�   �   �      2T  	�   <          3U  	�   �      �  4V      @        X2     �                    ��                                                       @   �   1�                   ��                                                      @   `   2�                   ��                                                          `   3�                   ��                                                          �   4�     �       �     ��    ��                                                �     `       �     ��                                                        �     �       �    
 ���   ��                                                � �����      �    	 ���   p�H                                                � D   �   <   �                  ����                                         <   �   D   �   <   �   D   �   3�    �   �����               	   ����                                         �����      �   � @   `   @   �     ��       
                                                � 0   �   @   �     ��    D�H                                                � @   �   @   �     ��                                                       �    �   �����     ��  � �H        	FIXED_ROT                                        �    �   4   �     ��                                                        � T   �   �   �     ��                                                       T   �   �   �   T   �   �   �   	[refname]       �  �	  l  �
      (   t   L   �     �  <    ��                                                       T   `   �   �   T   `   �   �   	[devname]        ����������������       �   (    01239:<      5=  >7?@;46    8 �  vcswitch     Miscellaneous      �?   9 
 �  X #�    ����11      PASA1�A�����#�   ����22      PASA2    ����#�   ����33      PASA3�����#�   ����44      PASA48 � ����Switches Generic              Ctrl1 �  b�     V+        ����V+����                        ���" 5 G  Ctrl1    Ctrl1 		�               V+g  	�          �  V-h   �  �         V1     �                   ��                                                           `   V+�                   ��                                                          �   V-�     �   �����                   ����                                         �����       �   �����       �   �    �   �����     ��    ��)                                                �     �       �     ��    ��`                                                �     �       �     ��    ��)                                                �     \       �     ��    p�Z                                                � �����   
   �    
 ��               	FIXED_ROT                                        � \   `   \   `     ��                                                      \   `   \   `   \   `   \   `           �  �  �  �                � 0   �   �   �     ��        	                                               0   �   �   �   0   �   �   �   [dc]       0  P  h  �          p   @   � 0   \   �   �    	 ��        
                                               0   \   �   �   0   \   �   �   	[refname]       0  �  �  T      ����t       J  KLNIMPQR      O    H �  Voltage Source    Voltage Source DINRoot      �?       ��     � ����        0      ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       �������� V+V- E+volt_sourcevolt_source   +0            E+Sources   Generic   V1V1          ����       �0            0      ���������0����      @5     ���������0            0     ���������0��� ����MbP?1m     ���������0��� ����MbP?1m     ���������0���{�G�zt?5m     ���������0 '�~j�t��?12m     ��������    �0            0      ���������0����      @5     ���������0����     ��@10k     ���������0            0     ���������0            0     ��������    �0            0      ���������0����      �?1     ���������0����      �?1     ���������0            0     ���������0����      �?1     ��������    �0            0      ���������0����      �?1     ���������0            0     ���������0 N  �����>2u     ���������0'  ���ư>1u     ���������0'  ���ư>1u     ��������    �  ���� 0 0      ��������                0      �������� ����       �������� ����       �������� ����  ��    �������� ����  ��    �������� ����  ��    �������� ����  ��    ��������               V #�    ����V+V+      PWR+AV+ � ����#�   ����V-V-      PWR-AV-NDDA����Sources Generic              n f v N r j J �� �& 8 � � � � !� !   L  � p l h t    � � ]� U � ��� � z W � ~ Q  Y � S Y| ) U; � � � W[2 . 2 �T �Z � *  ZP �  ): a� � y � {  � �< } � R � V �^� ( � � T� � � � \� X � XV                     
 �@ ����        ���������             0     ��������� ����      @5     ���������  ʚ;�������?.1     ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ���� true
     ��������� ����  false     ��������               
                  � ����        ��������� ����       ���������  ����       ���������@ ����       ���������@ ����       ��������               
                  � ����        ��������� ����       ���������@ ����       ���������  ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������               
                 � ����dec     ��������� ����     @�@1k     ��������� ����    ��.A1meg     ��������� ����       20     ��������� ���� true     ��������� ���� true     ��������� ���� true	     ��������� ����  false
     ��������               
                 �  ����        ���������  ����       ���������  ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����  	     ��������� ����  
     ��������               
                  	 � ����        ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������               
                 � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                    �             0      ���������  ��{�G�z�?20m     ��������� @B -C��6?0.1m     ��������� @B -C��6?0.1m     ��������� ���� True     ��������� ����  F     ��������� ���� true     ��������� ����  false     ��������               
                 � ����     @�@1K      ���������  ����       ���������  ����       ���������  ����       ��������               
         ��              �  ����        ��������              
                  �  ����        ��������              
                                  
                 �@ ����        ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ���� true	     ��������� ����  false
     ��������� ���� true     ��������� ����  false     ��������               
                 � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                        � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                 � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                 � ����       5      ��������� ����       5     ��������� ����       5     ��������� ����       5     ��������� ����       ��������� ����  	     ��������� ����  
     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ���������@ ����       ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����       ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������� ���� true     ��������� ����  false      ��������� ���� true!     ��������� ����  false"     ��������               
                 �@ ����        ���������@ ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����decade     ��������� ���� true     ��������� ���� true     ��������� ���� true     ��������� ����  false     ��������               
                 � ����        ��������� ����       ���������@ ����       ���������  ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������� ����       ��������               
                        � ����dec     ��������� ����     @�@1k     ��������� ����    ��.A1meg     ��������� ����       20     ��������� ����        0     ��������� ����        0     ��������� ���� true	     ��������� ���� true
     ��������� ����      I@50     ��������� ���� true     ��������� ����  false     ��������               
                         / � ���� x'     ���������     �-���q=1E-12     ��������� @B -C��6?1E-4     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x	     ��������� ���� x!     ��������� ����    �  500
     ��������� ���� x     ��������� ����    �  500     ��������� ���� x$     ��������� ���� x$     ��������� ���� x%     ��������� ���� x"     ���������  ���� x*     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x&     ��������� ���� x     ��������� ���� x     ��������� ���� x     ��������� ���� x+     ��������� ���� x,     ��������� ���� x-     ��������� ���� xg     ��������� ���� xf     ��������� ���� xd     ��������� ���� xe     ��������� ���� xh     ��������� ���� xj     ��������� ���� xi     ��������� ���� xk     ��������� ����    e��A1Gl     ���������             0�     ��������� ����      @5�     ��������� ����      @2.5�     ��������� ����      �?.5�     ��������� ����      @4.5�     ��������� 
   ��&�.>1n�     ��������� 
   ��&�.>1n�     ��������� 
   ��&�.>1n�     ��������� 
   ��&�.>1n�     ��������                 ��=                Ariald         $� �|p�|����m�|+j      $� �|p�|����m�|+j                   ����            �Fk               ��  TSignal                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                      	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CDCsweep       
 z{|}~����               
                       ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                       	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CACsweep        ��������               
                       ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                      	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  �� 
 CTranSweep       ��������               
                       ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                       	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CACdisto        �����               
                           ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                       	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
         )                 ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                       	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                           ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                       	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
         !                 ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                       	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
         �                 ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                       	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��        � ����        ��������� ����       ��������� ����       ��������� ����dec     ��������� ����       ��������               
                       	    ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                      	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CACnoise        ��������               
                    
    ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                      	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  �         �  ����        ���������  ����       ���������  ����       ��������� ����dec     ��������� ����       ��������� ����       ��������� ����  	     ��������� ����  
     ��������              
                        ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                      	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CFourier        ����               
         ��                   ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                      	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CACpz        	 ���������               
                       ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                      	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CDCtf         �����               
                       ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                      	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CDCsens         �����������               
                       ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                       	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j                  ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                      	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CShow         �              
                       ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                      	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CShowmod         �              
                       ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                      	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  �� 
 CLinearize        �  ����        ��������               
                       ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                      	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CParamTranSweep        �������������               
                       ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                      	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  �              ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                       	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CParamACSweep        =>?@ABCDEFGHI               
                       ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                      	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CMonteCarlo_op        ����������������������������               
                              ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                      	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CMonteCarlo_dc        �����������������������                
                       ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                       	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CMonteCarlo_ac        	
                
                       ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                      	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CMonteCarlo_tran        !"#$%&'()*+,-./0123456789:;<               
                       ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                       	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CACsens        JKLMNOPQRST               
                              ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                       	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j  ��  CNetworkAnalysis        UVWXYZ[\]^_               
                       ����            P               ��                        v(1)       ����                  ��                       v(2)       ����                  ��                       v(3)       ����                  ��                       i(v1)       ����                  ��                       	v(i1_vrl)       ����                      $� �|p�|����m�|+j      $� �|p�|����m�|+j                  ����            P                 >           ��   CDigSimResTemplate                ���       ����  ����:�0�yU>20.00n���   ����                       Arial����                       Arial����                       Arial  �   �  �                                ����  ���� ������       ����  ���� ������                 �               ����  �����       200������         0.000000e+000��    ��������      0.000000e+000��    ��������      0.000000e+000��    ��������   ����                       Arial����                       Arial����                       Arial����                       Arial      �       �         �     �   �  �  Circuit1                  ����  ��    ��������                                                                                                                                                                                                                                                                                                                         �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                       �  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    ��            D P��                H 4� �� . CE                 2         �  �              � � �           <c)P    ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                               �� 	 CTitleBox                                                      �  �                3�         �  @                  ���                                                  �  @  �     <   �  <     ��                                                        �     |   �  |     ��                                                        �     �   �  �     ��                                                        �     �   �  �     ��                                                        � �      �  4     ��                                                      �      �  4   �      �  4   [title]                                       � �   D   �  t     ��                                                      �   D   �  t   �   D   �  t   [description]                                       � `   �   h  �     ��                                                      `   �   h  �   `   �   h  �   [id]                                       � �   �   �  �     ��                                                      �   �   �  �   �   �   �  �   
[designer]                                       �      �   8    ��        	                                                   �   8       �   8  Date :       �    H  �                  � �     �  4   	 ��        
                                              �     �  4  �     �  4  [date]                                       �       t   8    
 ��                                                            t   8         t   8   Title :       �       �                  �    L   �   x     ��                                                         L   �   x      L   �   x   Description :       �  �  �  �                  �    �   �   �     ��                                                         �   �   �      �   �   �   ID :       �  �  �  P                  �    �   �   �     ��                                                         �   �   �      �   �   �   
Designer :       �  \  8                     uvwxyz{|}����          ~     	title box    Analog Misc      �?    9 
 <�     �  ����        ���������  ����       ���������  ����       ���������  ����       ���������  ����       ��������        9                                      ����F��� ����     H�            title                H�            description               H�            id               H�            designer               H�            date                           ����            `         �?�� 	 CGraphDoc�  ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                                                                                            2         �  �              � � �                   ����                       Arial����                       Arial                              ����  ����        0��          ����  ����        0��          ����  ����        0��          ����  ����        0��                                        �   ����                       Arial����                       Arial����                       Arial����                       Arial����                       Arial����                       Courier New                                    
cgs 76         47 80moh5.6 �@
KCTRLmvrd nmodel ATA
>DAT2
     ��                      TIME� # ) time                      ��                        i(v1)� < � i(v1)    TIME                 ��                        v(3)      v(3)    TIME                 ��                      	i(va_ix1)�   � 	i(va_ix1)    TIME                 ��                        v(ctrl1)      v(ctrl1)    TIME                 ��                        v(6)      v(6)    TIME                 ��                        v(ctrl2)      v(ctrl2)    TIME                 ��    (v(6)-v(3))                  	v(IV_VRL)� �   	v(IV_VRL)    TIME                           2         �  �           Time  � � �             A
>D    ����                       Arial����                       Arial                              ����  �����z�`?2.035181e-003��G�6      ����  �����z�`?2.035181e-003��G�6      ����  ����1��{��%�-1.075922e+001������      ����  ����1��{��%�-1.075922e+001������                                                                       �                      �                                                      �  �                                                                                                                                                                                                                                                                                                      �  �                                                                                                                                                                      �                      �                                                                                              �  �                                                                                                              �  �                                                                                      1m  0                            100   100                                                             1m  0                            100   100                                1m  0                            100   100                                1m  0                            100   100                                                 
                 1m  0                            100   100                                ��   CMiniPartPin    ����V+V+     PWR+V+g      ��   ����V-V-     PWR-V-h     voltage_sourcevoltage_source                          ��    ����11     PAS1S      ��   ����22     PAS2T     ��   ����33     PAS3U     ��   ����44     PAS4V     vcswitchvcswitch                                          ��    ����11     PAS1�      ��   ����22     PAS2�     BatteryBattery                          ��    ����R+R+     PASR+      ��   ����R-R-     PASR-     RR                          ��    ����GndGnd     GNDGnd}      GndGnd                  ��    ����M+M+     PASM+i      ��   ����M-M-     PASM-j     	voltmeter	voltmeter                          ��    ����M+M+     PASM+2      ��   ����M-M-     PASM-3     Ammeter2Ammeter2                          ��    ����11     PAS1S      ��   ����22     PAS2T     ��   ����33     PAS3U     ��   ����44     PAS4V     vcswitchvcswitch                                          ��    ����GndGnd     GNDGnd}      GndGnd                  ��    ����GndGnd     GNDGnd}      GndGnd                  ��    ����MM       ��������MarkerMarker                  ��    ����GndGnd     GNDGnd}      GndGnd                  ��    ����MM       ��������MarkerMarker                  ��    ����MM       ��������MarkerMarker                  ��    ����V+V+     PWR+V+g      ��   ����V-V-     PWR-V-h     voltage_sourcevoltage_source                          ��    ����MM       ��������MarkerMarker                  ��    ����GndGnd     GNDGnd}      GndGnd                  ��    ����11     PAS1S      ��   ����22     PAS2T     ��   ����33     PAS3U     ��   ����44     PAS4V     vcswitchvcswitch                                          ��    ����GndGnd     GNDGnd}      GndGnd                  ��    ����MM       ��������MarkerMarker                  ��    ����11     PAS1S      ��   ����22     PAS2T     ��   ����33     PAS3U     ��   ����44     PAS4V     vcswitchvcswitch                                          ��    ����MM       ��������MarkerMarker                  ��    ����GndGnd     GNDGnd}      GndGnd                                                                                                                                        
m1     8 8 mm l=100u w                        used                            �2�    �Q�R�XR��R�                        T�                                                                                                            (f    x=f � �'f                           �(f                            ,�e    �f � ��e                           ��e                                     �  � ���� �                         .I                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       h�    ���������                        ��                            1200    E-002
JV1.I                             G4                                                                                                                                                                                              �$�    h&��&��&� '�                        H)�                            MJ         W X Y [   Z                          DIN                            sist      resistor DIN                                                                                                                                       1200    E-002
JV1.I                             G4                              3 ��    CTRL1     
>ENDD                        -002    2 2 2 2 d                                                                                   